`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YIsgRh/j7ocOnaZ2oVEEl/TlVdoVauCGkaRXXNMRsNASniEPj5fyEqN6FPSfJT2QU8ebQqowfTT6
EFeDMujdEA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lcxbt7lzASoyrsaAxE7XP4Afm/Z81HnVTcc1r22MCXdJoXol1FUUr4ZnmclFBxxDkxjLIA3nwpKW
/rm9smYzcBR5gbwB8zNwGfrLQYWrBkfCoCXO5+YtZYGW0g/2LFSP3IC5wHTgunBjWH1WQqLAWesu
4ci28NDaoCz4uOLvyg8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dMu9sd7iRDJAohj9DNG9Ud+fDwkekxujClfVu2XRliD1ol0qPoVZU8SmFV6FlbOcRTll6IAPY3Uh
NOztCEHqU9rK/UeuTjZZ5SeczsGUWSZ8EQEX3YwcZw6gsdck2ljTzBwtIHLrD4nvE5xoNFx6XR1z
4CbzP1tZ6zpApHJp+4NGI2oCWZA+ySG3frdpxsK7Pp7QIt3Ncg3Iy4AdJEoE+bPdnptlTTC+u7YC
ladRP1D0/8H10ozzPfEMm9saA5KoCktpsBELRD+N/uAWboJaR+UvEgnEEsshDorX9JhPrNRgNjNC
ff8nW1OP+TrYbABqQg3RJrv/7a31N7RBg0JpUQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
vKZnWKdSf+vFEAiK/k4oUAp+ASSNUvfisKxN/xsWaJv4BqVAQxrslfFosgGOMaElEXxC6Q3LGv4X
ujWP7ibzr+NW/a1z5Iu87CiPzY3MfOgH6U9PVYwp18NsF74W29l9m+E3ijYfq1nlHktbLmoU5D+c
hcfJh6AZd9sSFClcbNk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mNuoO8r0k/T4a0BkWCnExUP+biIDpK43rSz3FAilgOmvRpcACd2SyaNOcN7AmId5p2cfnAOqCnux
NEM4IxP4yFvTDTEWAjRV1nM/zzNl9ovP374njRsCFq0adj16WNVzVTlJXyiOK4wPkbY0XDxPZjnC
cF42DLgrraV//avUqivs1VHpQGigGm8bYc9YK53xe3s1ZpN8AzaMyX6ycenvL+jPAUqtESpNtpBG
ht6W0h+GCo4+j0Wu1A8JkPPuMTe4C7iCF4r9szrbEPfweKpB2DQ0VKDryP5v6ogeFU/1TBbEPZQY
ss+H5e/uy29bSrb2aOv58IAMokI7jw4oZEktIw==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hUD7zFiXxoKCJOXjeKDAZM6zwXIY1BYdqxh/zdR+ph58scgMG3Plvo3j6JYUKzDsMeHyG5/FDR9+
bTFt6fiwbENM7XF+l0uJz02wEQC6o/8dgAvSkK5dmzwZE+zCSH//ir+aQvMeoVGZ3IdZ9yQ6x65Y
dvW767hyq6PGW0ZzNB4j6k5bzmwLEpvi37mfDHZeNhWZ/JK4h6brydPPGTYLXIgmL0HDbWm7p8uZ
DGxlcqBAe1m0aNcILYzKPPY2ASZoek7BtqdFq7PVemm3c8UgBCqkDJJ7avFCuEpfvAZPaDxmvUzG
eLYA5En9FTXZ2SucipcuqPlY471t3xv/W+2oWg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8912)
`protect data_block
JKR64Z5fJ7emmfNBwI81dkNTtngWjBSvz9UUBe6Ox/Si9VElxmCh3kznKmKkTBJVatYGpWUj28qp
FY/O4JQLd3zg4mnH7HyQHE3CMekK35fcig5Xd1x54sfLWCZTp/3J5y2opqAD7lWO5yTiVzLdVP+i
rIYB1f8mcZyBmNtg/vT9amiNuvbDqb+6SKe0U68/XNJ/uDTk5+wHJvVDGj9XearPCl65weiM2sCO
IsBc2/9QXuG3Hh6gcXIUr5JitABbBMQPUF/h5QrC28jf9sbB+/gMjvZerKHxCCADZj6IaES/2n41
LvodsO/6D6wlktUP/5hZ59Asq98qVvnO7UcWDwjKc/FF52afOfYFdgGmP4wCd+ZXDL8YFZPQQ/oV
S+GbrzoCTVO3Py9jfJXgYo6zx+sxSjbIu65qhP5pB98vlVvNu4Gn4wsMRuqbIBs1odSsdfLB0p5O
JyzW7Rt3svJJD3Llu9UPsd66svtT82TcnwOVpgB9rWtWObxvsBIPTrbXgl9NJruBaj+Z0E9Ejo28
fGwMqNTDZoGtLGDhsFCc6Ia3W07HUcyfrcHyf/JzQpeWUNypWeRHLT8wgjSTz5VyjnumQRhX4BV1
vGUYsD8AlSqso3wRpao9v4ZKyirmrCQIkCP7oN2WCO+uHZXyXxWQhuXr1gEjN+61C9MmERLe0Ksc
py6SVBKG0pZ/9MVFboNb3hX056+DAEw8RcVoJsY9+5J6MxSGMzdMZJpgZsHg271f1C0bYVdXwZY6
1SWJKr9BFdxjnj3zLcPQpzA147hWeObSTlEQDVdomQfACUYxprJ4jFaAp1ikH69Rz3VJ9BSjxqd5
otq78db0jdQ7UhmK+iKMt0t6w3KJn1WZO8FD86BrvjWIXL4q/F6eEN/KbklGdTW0X8ElyjAFgYif
/e7UaHlxUbhR3oRdgmbY+NMCK6vhX36ETyxA/e9jZiHxzsgKhzcawtwv60XIdnstkuhCtNwuQFav
n5BbGulGbHq0i8L8EY+mgVIHRyje97cpAJ012a9tEfDtCbuk8JRlsyG5ADIilgTFBbM5lqEQjw9Z
obqryZ59tT5ju97M+/pM33ubTIbxXVtq/2bflppTrFZPDfMkUf0xmeCPD7cZErScDdlwcvNQpNYl
kenAEUz+iBzg3FvbfqlZRN+xprCN1fB12a/8kJwg0hxUGrfi/F0eKJIPDAEdnSEss5XoM8BkEBu8
tbWDgGroRUCguG1I03Yfl+Mozr1GyTF1/2Giits7bMjpRAg6Enk1ahqYRpxFNXkNZeb2Q4nuOCaL
Yr4DYe2DKd8+YmheshouaQZqhMWEfnc3OR09c9bwSjNO/0MhhrhzCdNEJ99IfqJL3BkFaM9tDJti
B2kglXLVmNcc906ZdKNu86qYHFiC149fGUGHGH1MEX6A9UjrDkc7bBCuRsJ8v9EIxVRkzBbsTN/G
ZVhexziWQYljcU9M7GuD0yXtb4LvcxicEBcFkasCPahfOTO7ATFEOrOqd5NrEv89aH+p7qHRLEAx
6mCmfc2xpR79mQbgeyaR7wofv8RCdwqS+hY4Pw0Y/8OOX+FcKL8DDIpzliZhirrbQGuVW6xSesFi
pAver6BD2nSNQGjqZffFU3WZQepaGjCK6BZ7+t5wnN19e6cs2vbWZmJCwQCW0xcYl2Y9UYq1dVN1
s6h00diz4n18CLetqjE1JnLJ/c/qzGlG4vn2efORy9172oaz8zRCtIkbUbbK1o6zZDizF2zgiZzu
MQah3ejIn4M2XzNdqtT/7AeTZ5g0BriXsjXeEop5dOiQOZE3NBWDj59/uiRH2gyOilGbiiZFip+0
79bS96TrOjdP1pLSl/nX5+G4qnWc+9ti1KhSNSP+t1z9jd7r8O68LE6A4Rq6CwfxPM7tnegajj/v
hSlpHuJ3YBzn998hMgyGMu12C301moDhuCqtZLEh844cw52NZJ9ym7F0SFSMe0fJkPOPMtCE0+UD
sRX6cS4hleRWx6SRwFn1hyJpbObAgqCJOIkt/cpIEG8RQKVdYOrEPs8vj+E4xJq9tZK8trH/QjOO
JvH68b1POcgRP3kU2AagkMeOcLiFvkToCGkruXid25/19QrWbzLlwzeEnhVjJWYbTQg1lQ6csLPR
+YHaTFa/3HtjY3BJ5B4xUHKb+mO1AcYCd3tQmt29n+dL+YtC2lpMhnNriBbmP+qNNDS8nNsyLGLD
vD1Xr0xYihw7OvZjwFqwhAsWVQAV1LXzEKst1eGV+yEBQVCXR2rUSM5KC7GZDtTyYYts+htqlz3T
gv5ZKLQ3W3E+LTLgcEptHNZSWpoUkcbNT8PtPijGe1eQ8tcma1UKFJudTS1tTC4UnlBZ1mG5rOBc
VwrUkuO60fK78AxcExfR/0UVRJmNlvDSP0sYWNLYFFAVY5QlVnn6sy+ig0d3axIhi3ofylPVfjgU
Gl4YyamRnr7hKBWushP4BoUHJ4HI13HicbEZg8Sb+WFwfEpoePfv5mOdFngnV8AR0oVMnJ7XK3kb
k4srNYZcDRJFFmYCLc8MMgLDjfFQqe1VdjiPuMzWHcl4al/bxA1t1tjHotjHQvRrl8fhLV/0OiWF
1FaCE/FCtWxjnDEgvMgqYMh0e/AMp9tRlhSV1jM2ujL0Gp+wgKprZNseu8XRAogzf91EgwUf3d/h
S5ru+XxPTxOA8pRr0FlEwtjsvQB5seRJivprLDLlutyefg/+FKAzROyPqz8j2h84e1a4DBZv/4FD
oMn4ydHc23WPiUQtUz4o+IKfmd6S/buG2M8770KN5obTzw9+pDQJoev45GsPEFSJfnBVmfiMZwdO
bjbkk/b9kDlXRehaim06jcgLovCsVOcbFJbwLX7jBsVWu77ggBOP7ZvOOgWnykex7/mdBb+fVNCf
ZrVLqAw9kYCR9uQWOR7SY8/WLqiZcPOgplnu8vRvi2k3u8ozzpJ8tqiYUG1Zboi3XYQBarEmHk+S
YkvaaVbm8SK4X3Vvq5aolTxK/ORPaLYdARKDQ5xeBwE6wSrLtzi1ScXBoGO7xRkYc9/rqK3LlLzN
O70hwPJO04M0gzxfW89PsAr/AKZ798ssU+HPdTB+iGf+aqp2Do+tuYUbg5FjSgJbBos27AKaRz7U
fRyMHPsF9E+DT2Ae65mG35HqveEk4qB5al5GVRaDM5f56xzvf44jv7wt08b4RPQRK64dW842n2qR
yFEHgYwsPFJSfBShVmoxmkZfmxjiRn73yaUqEHhsmly/8uTsx8N6mzCkvg/OYcqHYaV8PrlAfNdm
rC5xFwYoCZcx2dBLvPO3kFhxEKpUYWvtpYaJPaell9maJg/6rZ1uXWmMwCCNkdeJeOrqeoydiP0R
c7HDcm/zjq8AB2MTZr5fNYu6Bd2oIGMSazd7S3gL0HfQlFf1lbUgu69nXM+ccjNKlQNsprFaWt2T
lav3vBYRHODZ9huXC26bTDHa8eGSAyF8Qfh5XDIrfQz8f1iEDWaFN+u09fhJ6v8Lj59uIiZuebkT
P5tcmgOAo20D9a0v2l+YpIEXZyggG/fKmLTz9800dpN3d1z5QDiMniG402wNlpHrZ9w1ZsBpqb8k
qfOm898JHynsk9FA2waw+59j1+twrXX3qSmazxZIw3OPAQ7t3Yu7O97qswIMG9easEP7mV9G2ZoK
3I3QmLyFBCznRs1fKjLZ4JTrEKpXHoewzqeXnOm+RRum6AlZrV7m//giwT3magv48+2E7JMcnuh4
hOU4Ei/wJEuyGYhGqVff8SvfGZzAXkbSU1hZvzi6cmL1vAl74B1afc8VhSfs246txv5SRvLBnv6o
5P8j+oxtTaCjckpzvypc/QFplLveTdwoMxqy2qG2+yI2g0/Tf6Q83nDNVEdsntwqiZnHji5DZbkT
6t+1JFLPYVMfpAkRpXy3sRHfMNt6oJF8UWMYOGUHH0pvmOY6vXM+TqhA/vSSy8EuMV/QQSkdSar5
Uv1MCdulJtesS1jzwtgx8OboY11FxJeYU82D3QxeX7P+dWgMCLEANWiaGvxKnioLsp4gIbGPqXYG
eowHNAocL56THCQ5Oh7IgmD3I4MMhzY5qspYpggkqqWnZOIzW8oMCvsYg//y0SJvRlnX+eKqdCsJ
22JVXABZa1O5bV7QtJP0A1KBW/bOBJtYkmCkFYcPQpyRsDs0DFikSKFI2gpS+e2lyoDDcEfagL1d
pMTVf47wY5TI7nqPhLlrQ0XWQ3qrC6BVdHN6O3PJc9N7949AYN33Joq6zMJtnfJhzL5GGx9Uaf0P
2usWZ+vqwcoCszw9nIyoSVV2z3LK6qqo00vwUpNqht9ASKlKEMltSjEYpVI0w2LP8vwOhspKeOEs
AfFl3Pn2eez9pVpKVG+iO0zJZoPjxEIIR/fRs4IPvnTFSj2TUTSAZiBqWW+bnElVkxI951rdMU33
aNfuTZrkUfc2MvqWNytA19LRUSBpvJiFphWgHybvHP4TMurgj3nhCFwZWeJpvyp8E2wPZlI0Qtho
ZF1XomPIbwjin0CUurAynM+d4rNipjlUgCBy6oQBuTGGmoc0J9NmYZ8pSgWZa0kbP6ytkBEDhkTr
Zit5Bgm7Y+wif/CzmtFmhUeG1ysPiMYwq8NPT40UMST8waA7NkbeEtFsg5A+B97J5/yb20DZvFWh
EqukPm6lw2DqT5oP47V5tSuvyOIN7zcBLMxIBvwpP/i8qaY3j1GVLAJTR0bIbFq+M3TEsSEQwMli
FoVNDQkbeb31szzQugEMP9wHgqKrvqjPMSMapltyLm49tIDHakW2LsUyxynMcusar/tZHaMOZQOy
wCfHmY30AGfYwXyCclCEsS88W6HO2q3h0zsArHditM2z/NiCY03/xzD+oliUOXbgTa/ZGrvBrEG5
KR37OzH2aYf8OwKOIyq9oXmcLPDyWdvaLWbk1C2+yueBzvdIbDUVcrB0uUCx+ZBlBgarb3Mf6NdD
7H7V6QHpSlBAg9WqCSL4XMxMaSICXoZt2miJC4QIvJmvSf/YBgQfs9wugO5pGjP+f8S07ZZkGRy5
OvsHW2cvcNjQLLLkN3MIa/3ISBO0Q3gV6oy/spsg3aEgyANYtkcOp2v5ICspQQiHnPd4HEws31Lo
GNRfaL3ZXVLsSYUTLSwoaJqOErgq16E0Vhg2hTEeHTbcryBXytXoXPgExSo/liFGDbgBtNLS7Mgc
QWQouL7bHoLBL00W4xqonpwp/k0CM7weVYWwL+ZVMy4vGm1NSjseNDiB5YO8g+XCMatJl2L40NYl
V6qfNH4WqmJ6AYCdKAxQTF2xklZ1pMn8ongEu6YJy+d0sa07M3w3SQufStuScLFx/l5dYnYms110
I2Hc0SRiI6DouGKzSqOam81Tfw102HH35p7OXYlljDs3AbcrpEBtq2ANxiGmuQB+N6UH36zn7Vll
6F/Jy05CeOn61MVQE511eVyLslkt3dNZ7ZGj/32pqPQVlVDGGHQi6eQPDYbfj7XjJazHZdc0QzGv
7sLRUAKJfzbbLGpjGZJYYSeCca3NWGGimMZD2lWzYJsY5B0Zv0AhCodf3nIulFJ4zYrqoqwUmRWo
53L6GWC3wJl9J+RcrSxnJo12iBzco4CJ7DcSutTJ1ATmSla5Y59h3N3SuEtx8Iy81n1fsr6JZuCU
LRG+iDXV1kfwkIPOhV5SC14gicMqGD8khPnKqwgL7s8UnKBhNT8CeJDsM5S4X6KSp9DVxPS/laVk
fHHQk6j6rLAgXF8Ei4jps94QLbwnLKuQeKpvwQyTtb+bQNdcXRoNIvaxXaR9S3eqN/B5B3k8BaKo
GmhRLqQafda31Dx06JQzzEQ9gSXuoPAy0+BNtgKdt8Cjs6HgVbGnPZeq+Tz/8o+IXQPy8EucvKH9
qxmFqUHZntIrEjMu5ldlwyWClrBzGY/kE9KNAVWWbG3cXV6OTZcIz22dIghHJNz2UNA7X0kLsMT7
bWsX0Itlh/jAzG+233iimJEWi0vQlo6DkTKmlgDYN0lanNzSxtk1ZDr8+UVIIjWEk++xPE+ZYa66
YyxIUh8pQsZ2YwH5hAKpokcdrWTn7K4q4u2taCD8a+P9F8TjAxdZRbHHB0EWVXnmWA4NKISWa8N5
6GaESv4li2yPgJP/8Var7jbwM/MZXoJsea9k1fLpMrQbj9gBgGloDFi+lHkvnwMVZeUD4GvKW2px
v7m6O3ulDi2TBPfI6B0Jii/mQRzSTcKEhYevTafcUIXnpyZxX9KqUUR9kx5XnjsLrL/KJXqbU6UZ
ASHlbB16lizcwEGTDCABLv/RtRRZZjsKu3HKVSmnq+3VWAsNs5DENWpAKuVNZLYni/ZYQpQQ+n19
UnPyWb7WRKkO7Zmz8CbrQfBfsrSUUBifGKif0zD/WyglL2J7osZU7dJqYj0TAEMmmf0AFvETul1N
5/l46GyMV3nq8DGGzCs+c7A7tpM1Y9HOhlbqKmssOG8MB3UygPX2BnbdBaSRsXni7PwI8G8k7IS4
zrCz4Z/+9qrQPGqvMTa8Cponq1fl58vNC6PkynVZI5wlD8s+9pCmHt7k4+EcucY7V6G7f6Oz4iML
yfKUsE0oiWoozf+QHwvK2WG1w1HqSv96qNqFuRKwf2nlEGScAXRxovIqblX5wxuLMe9a4cjrCrTB
qg/EfWlt6bJsOwmOprtuUicoTnAnkXGGlDehOE1UQKjCBmKdrkIKGx7Wk3iw9IFfRvK4B9COYJ7z
8Ykr8BoK9VYystXfy8N+pd9n3coeLkUBCHtY6778mF1/VBjg55QimSOHzJ0kwL/8NbsJKeoq0tCu
ctvmr0kO2Fhb9APdIKZbgR3fd0qIILDHljEAKoZ9o38pys2WdkzAT/ER2RBVzDSHz39SI7PUc6Of
RM9yCfkI0Tu6fEBV3ykYtwQH6qmzFD0bTC6qolXiO6xwZUxWotOHxXdw5zKkP79lhlpTU/rHkQ/6
V5F9axvdwzI59GblxIIyBkvaDCNDM9+NCq8t3ywiXewXjn6dk0RmtO5kfUTblS+W8iEJOvTJ0Upb
5BWqR//pwzVLIHrd9ZRRGbUudG6rubR+nJ+elrKShZKBsiXIT/Hywl9W3bBzVd9j0FhWU9/WjC73
Oe5ipZT31y6/x/278l7p4POsYgXTyYaO6+USL9Ospc0RmOVT519TxRMA/JDbd92tKWamKrysqF6i
LYOpwNovxpHTw7CtjS27FKg4FWj4nXam0frca19mGnXm3dm26nCm+CbNRLdOrA5yPfhsIa9x8omk
n65Ncl+/V/yZPj/qbSSOf+EEUCItGAiEsdmJHUsmEFzLUQ3EYq5dFS396afX8McPQX3QIse3GP5M
gRNFfG5t5N8IZKPOLeaJgAgKZS1WAmRHmuzMm37hAhmJAvBASxwtNCS5LD1TfwEl6VCjdNY7WjUc
9zPYkcPTuzPdA3tBTNvLsditrvM79J5E3gimnN2dAWGb9QSLQxzXhn/1qsamRPDgbDqr94DhNYab
Y2nkIML0og/WZh0gU1nhm4TqaXGV0tqRq4VpM/Vy1hcK7FQmBjJwlBbPo8DKIGcKZo81hwr00ql/
MBlOPQ/3dFFo1mKL55oZOnuVF5Y5m33Ss0isiI6CDxFNMyu4sy6AaXl5vAgg/QM4u3N0NCubDQaH
E3AZA6fFMY2m+P6sWtSSAAzHZ4QcekmtM3OBu04JkAMrMBuI5wn4h4trSIgaPLvTWnlzq7iaNnj4
s3TdVNM3WUir+7xnuVeB4ky+UXMNWXFFqhTs5aA6k3KrvpwkGqO6NUodk3lWc9LQbk9dJwyIVEFm
zLkro7mbIeyh4THEJ7mR+IekU3rNsmBbiSByPH/heVjAlInJ6ARudiS2EfO50thJmt0hXAHtJXbQ
Wr06W3iEMFkw1N1fOIcI0dwq6KaY6lWh8qb8g/iBL83GVyXGW0ydECYlLccMXHCbMndhrpAPtZIu
rXzIErlEehWijhpmNzzDcxxr5TN+fQp85GSXRwCyUgd6Lw4oBl6jsg4SPCNO7Xh0EoxIFzZ0/xYg
Z3pj9+U83u1c20giSUElf89eSUbQ4ZZY8/1k3AQJAVY39xAZGEiCn9hlItc4PONmPLfukql9ZaLZ
AKgTpmEZz/FkrIoUvFjOC+XFd+3sp4xvXiHcRgLokHoEJrjhgRLGQP/5ThxbdNAR1+fiQkCU+1NA
h8DiqwRFz57frQ7Pk+EUal7/L3FI+xeqD+4j1flSJhpbVNgtTvJttR+Noa9JQ0L3Hcf4etHxtNqh
X2BpBcRcSwxxTMrpQQ0nV1Qis1DKYc5TcJlSJeejGEqGh48zlZ10sNAlhaeUale5RxUk/B5EDPLZ
VfWbZKSkygiIuWqniIHHSzk5O9mxN2NbLzdkTzcACdDqbC6h+dUNFze2k66ln2KQj09Uwx+kPz+q
ltQAiHw6hl6w8l8U1Ar5mVAH7PnZaXUBbAquaGJeS8IWYh0SRyfWneFCIQZJE9jKVlzkv0mwMW4r
wWn8qBF8173TtLhWY5OQ5wmw0iY4ptQdh9A3AWsjYUSq4cqzZHB8aNfo0FdIcxEM72CWxhmr0+Po
lZJtA4NMuK+UeTVRfTiPi9opHVvXMcsYbURKpsWUXwfs9+4+GnfUhfhYX7A/uulYuN+amqsNE9jy
+fZ0HKDfvroFUjYYt+L2Mo7yCgObtSSjKcdIFIHtqxy+hvkA7CVXeM+dtmSvxeJqtyQNac5GCksN
WKDLilImCcIa3fjsfsjoWrfM1xCbkjBfx5Zj6E47YI1yL26fpOMCyuQWhyx93y6ZyogVzDfbDj8/
WUi3pnoicQCVeetoDu6sT8DrVXk344zyAOl5gMyaZHIn3hVmaKmUJ34ZCMfUYcTLTRvDs+ydyrNj
rmBAbze62fKfHAiTldEqumkFqAAKzoSLSj7AHfMy2QkRVt5iKAYQjS5b1mQtqv1+I8I1itlldc3Z
uVDtS15/lyp3ZObbZAhp5vc3RrEvQOvzg9zSr0ZJeA4RUCoTqaUtbiy9W5yqQU4Kei4T85BcXRG+
vw31SMeVpD0Pyq6N3+5oIcIE53fpgOTw33GCR5g72PG54rOfGZ7r7vv4CDKgZ0UJntRc3doq5gNF
Jc3QoVWXdZzExyv5aQFq+Mb0S2TFg72BT+WWwuig/8DX0Kj4YJqvTtDVwM7sQ/vLM3gQxqC7lCJL
2FYwMCJUTeRfhICpp393hVdCeRPthjUjO4NbiszZjG7pZaZLfRP/80sNI0S7hR+qo6OtleZ+dxtq
HFRk4qCGvSRvN3vcou5B+Vb7na9jIiq8xrEN2CfMU4KuJaTNk0w9Zz511ZpRtH7eJiBJBJPa/cEW
HHN8l3jSqsm3L9MD/PZ4VbBFNSnyzS3n+/w+R0DUZjOhmmg6feHUf9C/6LdWF83/yo1atbSfPyEU
/gJqeDvBVBN9UjwKUeiDDGyVXZzm30Q9lo5yby5T0GYprh6OT6M+Tvi+vtLg4RWxkEu3HmPIiqR/
dig+/Ux08vGuBJdWZHa+iv5MiDjqKTmAuUdUF4eugiq+mJ3oC1eD/4N9qD5SxHSLTXWQgpBfJ3Dj
7EHJXAw3UHumN7FXK2EweOEcXwxo/wRlPc3ZHA/EFpxkIPetJPfdAmx77VsGJB9GbpkfbHMIvXVu
Efi6/4LfxuTjxcIEncdBd2/n/sWtt5Z2me2XFyJSXhB1kC2aXrWRHRJAlW8oAx6JHKXlIeQMUY2m
AOACXQxWrygKiepPiwUluWAfuGyoNH86HMHO+NWVQLz5jN6VNV0aipvmMvOESpVloefDBCFzD0o4
LZ5d/Qb6homyUJb0oKhFYzoZAfBU8p7XrsJS4r5GDurpoc/PQnI3sTg/HgXI5ajhLqKHaYfBQ2uJ
NN3NLG6hXvoz+gRkkuXY/+5+McUtFgCX9zV7m3UPGKPxEe6EhxsrhqTn6FrMjq9EC/R03dsEFpyH
nkHJ3fxVk4+nrCOqXrH82RFg6JyYhzGiMQQqb4irtyg2mRa6G6aGUs/cyn4soQ8qtIGTx7wN4x4+
nm0MPpfiCU+4hU+sxnN0rFXuvSQ9ZN6P8hz03yk635eEZuYGjE9m5aYqaeofPHoPCotHkEJXnWS0
xs1ek/Xgie29fahbHjdHaBujte0sToVXIB3YRKZapbF4vLvZwX/hfxs+UMBaTGp90kc5eCQlPdzT
pr7zFsqH8UzO4Tb/rRhLNs/7G3L64rAjS5LmZvZl+0GQIjXydNm2vHAgf+2z5WTAzgEAnVNJGLwt
ZaI6//RQHaHFEmakT2aUZna78rRZtV0BKaKhkwL3JgBhlJE3tFMD26b2uIitUj/2gAX+s39cH1Ug
wkYQlgSd/4KQvS+8ASIsy5JazwFMKRO5wknhNP8GXps93JQs1Km5j8wXbIgKOOr1sTSx2C1kfqJh
/OIlNZMz5v7Dxv7v1ItEaZmyqjSj2pMeF1cYcBhb3LMQ4reO6jnjPBQlESnufK9KX3Z9upP9IxOo
lbsrud+3oRjlARYxgZKtOI+ITsBjopSynXiie86+cb3iH1B9OhHufMNLElEljJXng/9ZlMOgK65T
Pmqj/JdeJZBJ8ZbGcUKmsLG9W/KUZ7YceOmCnBaDtbdw9+D38yKHr1QdFroBnguBeiWHYECpdVRg
f0fhVIr+F+VhvLwdv8mEEwstgJo9m1IaENkXmuBpof1xpTTyFHCv5CB8aPWz+TVgXX9+qbAJvUrm
Agpl5yGo51rs5Wwuevxl5JniAZK0fEpV9Bzr8qY1D6LvXiYesTa+90OMo31HXK8B31zjFJSXnVOV
lnh9K/YcFFzvAU3MoekbexIZO7rVVN0KMlUomp6mt1PcSVV2vsFGcgMokd7fLWurHCBnf7dFikGe
2/FKCtI+mcVPt6h1qXYQhrrYc0SkgSw//7vk1ThIJNf4/2d58VwDNnSnTiimI1q9Ui0h3TO8XTW/
Hsvl6emCn6cfv/CVN38DzMCr7QPBhZi2U8a+2WAw5F/MyXp9eEXvtpiI+qX4rJ6fV9lFlefadX4q
DPH1bo61HTtaFE9YbkEocCU8iGx0mpcDizhkkCIFIU+jqD8e6RpjmbqqrTkrbzdYfob7yvEH6dbq
ufLMFYr1WzdWBBIx2RaedizofCWa7u3sWVI5fKtFRpXUChu2JQ/vpumeES+YbSm3oNT5pbjXpDlx
1S7jy43gWF4SfQbBB42OqUW0yFsARmNV6xZcjKT+P5b16M5+uJ89/akYt/VbuSYMKipoXHzRZL4T
k5dhuu9Gg8B6HHWZ+eRobdVtHP47dSubUBCvm6+z6kczeoMtOPuD7pkg15LEng49B3yEd8r6pqOp
sLbAYcxpeZyLvVxfX9NRKh7OGD3AnP31XFdzgdFwSU+Cte5dNhOYTUnZFS/79N+U0luvo6Ohwxh9
KgW8rZrvR33kzCPwV0nFbQj6pRFLkdV3OpnuxwjtUJ2f1QBsiD+oMXCAhM32b3cO8Lb+/W50AN5a
neaQduyiz2rlG0zMEmmzpqROSrLAt8DnwyM3vesT+C8luMucoKrxNo5HTLQZUAqf+FKVxP6Jpvgi
T+X7QMVgbwqVKNINguCGxExU6GyyhWW0hMkmc5I2jj1hVNS0cROmTkiZloSY4lglsaRvkWcwrnXM
CE+rN6iUu5rST+30rqTyaEg1n12duqfNvxgg9YY8/uGjVFk0DGRpQYBv9k6Oxqf14ivmoon+2ZuE
SePcnI96sui2S9JBYXDdNIwBt7tXFaFX6OANJuJf4jQ9+ke3+1dsVP8GtWAn+kONJHLhRTQN/445
dm0Y1oBU0SSKXjXnl0uQBJEgpZ3IGYkikn8IlUxkJ8bWmqJ3to9Xf9O2tM0o90fYNc7n+3Q6aZnU
viAW0vLGvItaUOBeL9GT3oA1yMJMBadi9Y3wneIn7HS0NsalPCeX7MVW6/K0PZyn/8vk6HTVXctZ
m5xW4QJyD85U9UW+p1R98a+SOgo=
`protect end_protected
