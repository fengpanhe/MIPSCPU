`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
T00IF1U62zm90btmtEJP5pUDXdT1ffoo0sDkNgV2v8Ii40nNNBuOC9K1FTtvFetqPupcEX/VGFR2
MIAViadEfA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
U+bSe3zRBcz3iVkQlIia8k9wmbi7gWNt3le0vDSNQz9iU3a4fDadlqSLshEumal1ic/lvogn1xJH
yTTamdZrkcE/uG7a1+2NhhQNKUj/ZG857rV6Z6v+rgJZcnpCIeskcbrAKP04hyviOVcQnirGPP2H
YkjlVO/pyYYCZnuQk7k=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
adqdcx+NHQ0j58sflTcj/3jLRM0rlkBvx+O3wLFiOXhiEkrsD3qT2LWL6htyyIpRMLWeUS1rBx8U
9+iyzsLMox3ueXBq5sgXU6eAsPyfEzH1Il9dHa/Bp4BAIVRrmsmqBVKry0A+5Vlt1R2hLX+iQ5AD
k5vNvxU7UEr9+LORDrb97j+W39z7J+Avhv5JVE4Hru/hEL4CQHYFs/jw0e+8DrgBmL8pAwmAJSH2
fk+0QFu+ZOiMeIUl7v/mntjFKBuauDorZFnRKOTOEN+ijUvY4FIm6/p2PmZjL4LIlp/qWKdin+q/
ziWsvIwr+KtA/vagPk7BqhqldpeG32XYuH811A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dxLiwmlgoL/B9W31QiW8HnbPOUeguVZHpV3tRXP4USEbanh+6W3k1lpeBWLPGdRC073CtoSc98b7
Xdcd0fy/1VDnOjLZHAg/hT3Vkb5HvbhuDvfbtbzAdeMbUKctjum+jMpyv5Tgiw0Ng1eiDAlJr3mc
2e3gqQ8ZjJdgIrqiI8U=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BJif77ziF7n7HDXu9iYbJ3bFFcDmf0eXkVftjuNlgk2upevPEcTsPHy0y35xv3U08CcBsTvD1hzh
+ZlZUjS3WDdHraxIbxgZnO82E1nRit2PvL/kRaGF5k7b/ZRLQIc9V1sLLs14Z9QNWHqrTkfCnGUh
j9kgJbBjdod5qYAvTFcuQDHY+FBvNqqNnNfTV/oTo2W1wUL8UtVhuSukhtzFR99fZguPWx0oPpvs
cZa8R2C9DTSPBKyZNaDAZsrF0hj+l3uJ+PWgKJ6LjR+azrqRH2vbZ04F50QcSYNZuevlFRFlHISv
Zvg2tS3ZSJCaH9qE5f9UBHsTbbbtEj8uGAv3VQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
e8T8l1agdAU8xGmSAUBmV+/OKiYvSlVX3Sppk3l4ZrWCd6qAo7xmiMn80RORrljpuAQY5V0IKVY4
SUZvG7DMuVHL9thJQgfSS35IzRpR0iN+ZvROcMC42OZJ99eJ7KG2zTMAM6P7w2ukTaRQf+UF5rpn
P/Ck7g/NB4RdAon9RKHlsyk5d60/rGLbDiWvizULsosxcrU0QOyKAGqA+GjNuT0iNsI6xnPQOCYP
BKvhU3PKqqCl64cv5KtGfi+e/sir/Jalvb9dYQWeYEE4dYbc9ZGooypgst989eVCwZ7lBVR/riW7
1fpvUTttxWbeIZEKq5S4/A0sUyNl2IX6O8NqNA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 57296)
`protect data_block
lUxDJVIwuFIPQKO/I6E+8DN+vwK/K26NYVfMV/PAijUDxEcTCD0BX5mwzUB3m85WtLJm/5An4QJD
9wMRlNAg+EQPwW721hdex9XTg5up/tTjvArc+37dRMraQMVskim9LxtQRYO3E3Vc/1TUSGGEX53Y
463l9OTaZME2d/W0lU2qr3o+/EdASutwHttk0vSSkzPrkcMWBRqRk/+P8WKyi6jNl0MY4qk4T1PR
rsefr9FLba4DRLU4Snkq1gU8KceBq1OAdM+qg64L5gTo9Xx6b9jCFI4+Zet7d075YD2DBhMfs2kl
038+0Nn/5Csv9S2ixM13owfms0xwehHRotQLswdHonzUzjspbOlMI/ZytR5UAiiltN8q1AW7KUEc
1G8uC/phyPizDgPhjjR+7v6DUoonx298kodiX1GDMzMRoZXoCV5UmdziXRHk+4xT/Aq3wwDUbeJQ
ROhkM+/s3wxGhrxjQxjUYnRP6DaXDAP5660zrPdiHb25UG+bJkclPjhVLMfXXaLG+XI8OmWGIZ2e
5aZRybPAOMcOoLmt/OrOLCFzpIhznyRZC+k9fbeJafBD/i22jU2PBVWqtb/QVVaFbeHGSSUhMvPB
ea/v9lXRINLocE5sdC5qwKHvWIQ/lBynHy8B+/CIu1qtrrCxPbTDSnOAODZSAUSWo3+YJfV5Biax
dYTtJrt9M5Yg0BzE0msfxNxmjK1Cp5lRYK//V3xux0R8bMThBrWQPYPh7lO8RDuwmzZVWzkrQw/b
7cKEbVOg6NAUeX5qd6MeZrHVvOmUvZha/VtyOqZ1JG6/UB7GjbYoBjIXNWKsf/DEZl4AzRG1xzJv
7oETpnWaC5YNt8a8WaLmqgh/HMsq/DThUTDeQoLgiQG47DUZG08tbttWR3rVtkLd4zI5ibuTzVuG
Rz92KsD9lcL6LX0qr4jt0ooltV7jxVmzuSZ9w46kAOTxGC/4IH7DrPSSRUnQeISMF6p2ff7H6I9C
gcfQZ20Z8fzAMhb687SSrYApB9aOjDTeaVTUOuMIF+mfGKRgJnjeNi16YCSSQTXDWnCOcsvYKyfL
ut0LCxKxPob7yMS3jK4YT7JWvzXmEO4upsG3REBHO0Fznm9b8fd+khfF01QcrNU965m6rtzJNzbA
6fAtw2Om47arpmedSh2pMybbSvwWk5HTL9aySztzHqxZXVGexvp1zerHvo2FqxPTkm2cPTFnAWnq
yW+RD2KOrCAnhMNtEcJExY8CjQI2amghe/UbxG41AN6g6IAqisPanM8USw9l1ZwoxWY6IZ0BmmeI
zXtSkr+U5vh5vTDKFq6aXly30fv2KNSoYuuFZJofoo+JYZZnHHMnGMWSIBm4FApZO0Hih+EuzqRs
W5oN6pNgsfzIDz1luw2Fu7DXtwvVfywHEf9SuIkJbq8qdirsYa4ESGZOcX6efnUYouajET5gUOqc
347v93D88mXPMmYSlEAMBHv5XNvZGaPshpPScPrc3XiZgT8O0HdsMksVaJEm+t7hZRtuxTC2Qiw7
vibl9IWQYub+fw+/OQG1gmKvmrHgoqaP19LtPt4c1l+0u5GhudyeuxZnmEUQi19R6DiehW3gdsOE
dO9hZBeTIxtgW0MmpG9Nif975hlmtkmDQK15EDq1Tv9xvISvdlYUNRIlgIDmDBaLI87mjgRWNvHw
coRGup+VvqGx+As4mOjL8RXd7Y8B+Eezci1SkeR9/aiLdwj8mbt+rej06B5Y+P0JQMKW+M++K/Qj
AOJPa5JY3xouy1t40hfqjucspPqDnKYLfhXPvXMDF7AEyMGxQB3qbLCRcuIhBOBrn7PYe29OJwbC
7ycKPOsUgBMgLW71qMx3qBbIfUhefgxbBMPKLYOkHln1turlC/tMePhhfDO3PI/EPmqgqA8st3d7
FDP7CqEDVGVhuM5Z3/M5hbNf1ehOqMDej7RWoeRvXEMsf54vLhtfPBD/wljpWweKTKcQReJk/ssr
vhsDizxF6LZUtRB5PiGHYcfeSml8r+JDcjnflE8d39GvVxsSsznUxfMhePiYKGGB5v+fyByzCSv3
UZZ4JHtPRcjZNaRHNNFq5RiW41e56EnZ5TcrqW1WjJUHroMWlOsyulr/g/aDTKTTcSdtA4cCyAmM
rheZwtvPM5ywo976gq28Xm1n3v9LtrRvnlhJahRXtcmZcr2PX/vayEqYuXU3RZqHNEpUCoNaoAEa
Ys5p0cDR7DgYjy0WtftD4Hq4SQIL+ZbkGT1zO9JhjbTCFqrMuB5M5l+BRWH26UgYuBrgFcvmMd08
iwrxh4hPiZYfE6/GldIswP6z+DWqX7GWX+RTU8yZW2tW9cxB0xuiebJq28wGKuvSlX768sa2EBfZ
v9pCcbeoAbZ46zK00V3pDMHwyFm1hDYyq8LfkjFcquHuWIjr0iaU9nC3LvgioqSdoVNXmaKOpXJ/
k93K8Hy7AhDSgFWdGxtIgrchWyuHmrn0uQCqhUJcYF3+cKbWLvZMa+G40OoGmrCqEUISTx99Cm9s
8aoMsCfOZscjv4J+TAX+iskO03ECHgQ4efPmxIWQVPWv/OoaoVw0VRISYBpnHBpQCz+gzI3soC1N
zRHLTUx8c6jebOiFVX6etp8P62Zrz/kfsjCu8TBNFdncOPZH/59W3NtQlvPTp7ol/az5th7nP8qD
DsmJD8cImZyDyT0qey/hw+oUKEQs6IWXGn4cVJRJj5CMnpoBXzwlMX6Q9Jq//vi5S0LHSWZWobEq
L8/dmp85cC8sNjg8UGeHBou8YqDEC1ug1H6yWpxBULPvuytgur+s1yBK3NNPzckGY/uscuQkQRgh
qPsDq4NGoaPpUxO6RCGxuU8l/efpThkADp+6N2NqYFXBAEKpLL0x+H0VCmThFM98xkzPSwI5SoF/
7xPw7wZ07akFntb8rS/+Uu1KenDnHRc4Ovgjh2UIAPUjbVsbQN+zf4Yj3S2FMtFG2clUuZ6SGS8f
v06Py3ezxPW8b02utpZt41wdWeclLn0nk/VNv9Sba6k2epYAvSYkSUuf7TyPCxHf0fvIr85kkx1L
WOWF0BPbW8Cttw8CHAuakIctM68VZxC2LIKpH+bMmcFOQAE9hUarAKlTjA+TGSOkJZNVzUBM/BD9
OxPlEXNiD3ZmK0swT4sniTw17cYN+GEWIS/kNcgDyotKOLPE8GEThgggX3RvlFxm8ETZsIJ/Xxmi
8CbtHju6QohXrVfB5i0JxNTFsxhjkztInRvMl12h7PyzzZdoHOijQowlfoXlez6ggQgdm7v3kQV7
zZ6RV6dW6wjKQt7lfBYNnES5PhPEH3vpQ7ZR+tSvnkhWprxRqs2lpDQzIk4ulQeoBvMaVLKEAppA
mb8jE6ywHCn3KHZJ+EcOT7P8ry1RzXLUEmHjhWVwZf7Ho9FsoCVDdy2WMH4hVY6DeiWZinie60v3
2lYoadgMejtRuw1WSfePhu6GpoiBWpSoKPqwYBPh9vo6tZ9tFOcsz2pcJgYXHhuOG7elraIWF9xe
TIQMJFaCz5bwxIXeFFyeqSfaFOYRwgnuFIDko24PkY3RZXWQ3IjgKxmuqsnhFB29a/CIo98zlvqj
27tDv/Ao/fhc/7a5tkdbyR2bnf0v5dgWBAeSUD748boFfLqfZIwShiHgkXeSdUYCev+OJVZnrqSb
B9Syj6FybkOImE74/egC2tGjwuvYHj1CY6GMDlHxmnPrwd45ucNmpvuFt39HsFwfGdt/ksU/HrHN
fP0IxCWG5byJOBuGRg1017G7nyXv2DwdxKrLNDDfBba8QAlFovhRzLVpYROuzXUqxTpTiUSSl3Cy
Hd19l3XXCohQP9xdb9veLMRcPXyNlaEyik4lpQ7ovUCkiC2yb5TFcHOhOgqbYVvtgNHm24IAdIZj
At802HGXMu7mdEeErMHXpuSSqaOReupTZBbijhaF/Nq9gqs4K+fostkBLeoAm9v2oRd3HW5uBXSF
ZoIiB5U7Nr3EHQUlFF2nuTOHmFYVSh/EOLF4Yq44ChKU8tYeBzA5/Zc/+dHiuAjFPkQmi7X/i6yJ
2/mCb0MUi9nsle+3xVMC7GCHGaepA/sCxRRFrWl5bN+Xec5kAjD5LKhXb1rEVDCLJODMgl9LsCu/
viuW1CJTyWEJLMJLbnLT84iagPN1TJVRlUhkCWqtaDE5qaK6D3vWu6La71NmnXw2JINx0hO4Fl55
C3ylCpSEXkWR6Q+mLTU1y4hlUb1fWgUGG6x/u97uGidCbd4RhohhUtXgBYSNYIo2HYute1edm5YR
9CNDoTvVAGQxe6XgpJKW1qG/zyEyp+gxl5BVNv9e+VpDpphCjkJt/aVnVUsU0KdXJkZJaCGW1DWe
+jHrf3gXXGYhZYv/9Y+LW/oSBbjcHqHCG/Wq5F+mtYqfkjaDOQBOD+in917XazbWJx0+Z3tLLkVM
ERMDc9Qj1/cyrOK9SGZ0uBQO4+OOPKVa58I0ITZYYMvRTKxdVjYzJB/i+D9ZiJ4YrRJ2Y63jSMcc
RIzM4X8EM/FjptC36ZxrMyXIcijMomwUei1jwemdv8H1F7h71ZQT2hGmiwHIyvRvJu3t/MTkb3y6
npNPyGdSueViETgSVmHlcqkEu3vB5LBYwf1kxxgdvlLJnZgoG4TIi5YqiIBCEKOr8UTmJ8WX/TQE
t6olRbxlYLp7wtpwVwmEIttUYwzuRRW5dTnPuomX7Y0aeus+qjFgy6ljjNsFJBMJ54nrcltHHEy9
gLtJ1iJJyI6BHjX4kHVffUlWSVsoI7Q4JMJTsM9pBbpVUBX/7Oj/z0ChyX15ZX+p4sVfVzXGA/sH
Nr+rxfSugzOMod0Fv9Tf6xmruqFYMIStTQxaYnHBpbGHEXD3/ysVRyQwz8HKyFe2EakrpSChwjRR
PM+nCUCN6qroHbHW23gSOr/0Ng56mqrwVSy1ODIQsLP0MIy/VDds0ltTlPa5pznI8esRc8uiWYE6
PoBNUNLeN4mzSDHslInZ0foXCbpH8Fl8YCCgBgn7WaDV7nFzwS46GjHz1us04T7s4XO+v30LigjB
ZRQjx4Kn5vpgy4D1BNdUu0i8Aamp7mvhvyXQugjpnYXknQmkfuHHAUoiOMb9vIww5RFeX50a7J4M
6pLQ4gc2F+s221eqAlrorB2VZyTrFCd0pYTXcsH+60PgBS6ocZ9TLX0BALQlzl+uXoErevPX78vN
P7XZwTXaApJu1P8gbj8TJKutteB//cbYX+J4PBwZIF45YlVscTPTcr/F16TzqEWK+3tPA0H9rcPm
S/12kkVyrOFkK0wliJevjPqXh70scIF3hLsOPR3LWF89TP3o2KvY1eeGGd9vK2bShwR//XKKvcVl
Swb6lQDxYFLWXIQhtAbjLLI/oWbpmwQ4XCdHDsMbMZaQbJIrpdxvs2ygDfLitfx1WJYjUa6xsKpg
yDsTOlYc8zOqV+lR96t8lpcpc1QsOhfglRLUscv4YmgNhS3oZlInpk54KGiCdP2iZYcEQ8ewFGiy
iUSS6uhcbAvrnPOk6Ql9YiaAP7qgCRGE5k3pLkuvbcorwK1WddOnArE5eJfPbt/6rkWSnftjfnYO
MztVH/xPmGY0H0qQfUBJisMYT+Ig1xCqjbQQJaUlCp46j6x3XdiUfxA+JfERt0CNj9B70V4rYUB4
PH1nEGj+jzlyuFNvLbK/5pf6DJpjLtM4R3FlRap6ZH8KeBsRvsnIxJppdkmxnu9s3cW/p5oLfU8N
/MdF8sWZJuV2jq6nNFZ5MPD04KWFoQhId/cAoBZTGeE0jMmmTSvc+HUb7X3MIVWIryljmLSWl2Dz
n8KYXxbrmwuHT7Zd1aSwZiwDAoom7vpy2KLqd7SWTbH1M9zkLH2ltYrlWwkOlpuzzOYvVko2/klq
FBJsYDq1XpMmXs3eHmIUX3X6rkCOK+h6CK0N1zhnIrRoAcikt4sBOG7svgwRDyd8pLC09oCcSPtE
4PVNykMLNkvn3mKiKBNYc7Enuj87Om25u1Zo/iZn60giL1C4ouxBJthoSmug4ciwiBgkSCcszOQT
4W6IvycSVVPVY3xun/UrqzwbSakI5fOsQ6BPGAfXidJiNzGhU7kKS4BBGmyUNIceFfzvW4Yxk/7r
5KpHeOWur/udKBF5fJHO/VEqyMxkUeY9jjKk5U+R1T190xtl1DgjYIN5yRATw5QkcYwG9hDykXIt
ZhLC/OnXFDKAef7YHFltIM2PElCE7sKC/K2xPKsvxZFkaW6l+7Ww62aZ0TYkeOtCqYpC3zn016eS
yTBU6x5V2N4TNDHmzNCGo1NMr2P5E9+P55QoP424laH8ebGd2+RFlVoiSyP0bj6L3ZATkpLLVQnI
3XKkvT8M8G+OVnGMxV7X+jQbRbIreCmFStt/pWxZ5mlUoNYEtKovb+xZ9sCH8/5mVa6Y5irhqXKC
0ZhZjFRMMRL63WJH7zx3LkjkbbPxzFA1b0JQL0A/i9ZPQQRz10c4NuKezfyZROVuzhSrPn7RPgnu
URdMZDh0Cbhrfwh4UQyJntHEe+37fNMDoZXCqcm8gXeyJSULy5y5fCqX+ADzHx2B2/27p1Lqbscr
NFjONDsxpvA/iIOwee5EB7DFXFnEfUzYYRI4WShsKU+/r2/ZszJxc+JVAj1oEFRcIcVVtBA6fenl
ruIMraD2gQxYwlo5EU0rhYMZz7k3abnGulV70JTPZW6sp4h4GeDNz6pNilOYO97eUxAOfTB0fimI
bDof3mRq89zTYbPfhz4xncuxggI/A4h1ZqAakuyFnCkK0JwAWBh35S0wyLh00nJ73OIvQfYhwy7c
FBCwE1oDP3Lr6PjpMxjCLVr+bLWO3xOiqViOUMPkmWKbWoIA8cZeeoFEd5cc2ye0w2636sW+Qbbt
rw5XrlfBjLlglpYykrW9Riq0T5JYK6709/DTI6C/wgwQFTDgkqUS0pJnpp4W5FzJrghqYZbbOzgM
VZarklRUJzH9+T0jZVs5SgtFM8LimzLvxCh0h46bCOrC+YrPq46IG+9mxPtS3UElQ+6UJ2c7WZ9i
24L5s7ifXY/od9mQeFBgyJDdWbOq9a4J0a1Z6cfKo1Rmn1O6Udyl/7JM8Kxg7o8JkpmPrT3oo+tL
OmkJyG2/p6Nwcp6+rAagS3vPX7gGg1e5OWA7p0sd/o5mURWLc6RYopOYysdaZg/RwPostjDNxZQ3
VHZoSDIl45Vft/Ifks0uboknFpREEkjr6Pl7JX8rNMkdpVAVcqRXu+2Lw5x4TquMRHgHbfGGTHTh
OaiOIvsMdmf6LzxPlqa15sK7PQqT9CgrcWoVjLzrjDReEDs9e08HGMXxsgiokic3hSUVeayQ6X1e
0CSAWbLg1IGxVDk2kZ109JTxn3uGYf9DpVt/3+cq1q3QWJGSSJRehWo6SyLUlUkfr9/jAtO4DqJV
xcijKcgUsMWts/ajYkVArFug/mBueIHqbOo1RiGrAY3WbJKp+IiTXD8mHmrGtmv+o0zK3fSwlF+R
DQMyH6CUvwGKFxIcjTO+TFHclTyN5Nrwz5nLY/zqtIxv/uEfoDLhRHRV6jt9hOwtod2ClCbc6786
AigkvO/d+sXq6L83vygyWix06x3leqO0w4i3PIYhRnMkHWF4H2/wDXhx8Pzy5BgaDk1XD82F3ku4
7vzuj7nG+Eavuem39fRh/LY4LeiMQ0pT43XfD7ATMf5hbbDgqjo9L5q9dSpwnpd8UqA6fSjxStER
TwbXb8+72+XbH5Fe65hp0WxNsqPD6D5CwAMidIzg0vO+E0oai9fdkzoj4lHUq6zMJUJWlC2FE93+
DzBziRXfclfj2if0YwD0je05/QlbZnygtyxagsly4H2xDUXMvtFVEaFuRpc/O72RJQ9nc2QtFNXA
MBFf1EuUJiS7A0QX99BnLHKiMLQQs0hN6XqO30jr4jOrJn0M+NK1oT9qcCZJCCpE8o4wZYkH5XSP
0pZbVr7AO4Dg8/QJQOIVR3ZiE/2bAJm98mc3sF1SIheC1XVjk7d7gp3bp9fhMdrd3hvwzj2SjZz9
o0zLaSjRr71TxxUKEaEPC+ciaKgIvdXUsi1B9KHL9MaFJhQIruFwFgAcUwuLD5S/uo9qqdpc4+Ot
jzxwwLtpZAI4tFNnQU1mUTyI5wRK0DY2DBZ0hCTKzEYO/QvvFASwXaYcJ5eCieyFcOulI6WNKWZ9
FN6nsvBbFR7334rTJXHOajIGCoUDd1qAngVZIb4WYulPzrLnfPfCmpnLCk5ANYmPrajMnrigX8Pk
jKl1k3U/2zQsCD5ynm3BzrbIGB0jsrAcqZHc0mRAEe1siGtyaQZqNP71GzQTHE/SZ5uoz9Y7YYfS
GfDS1qAF2sNjyU39HwTSgRK7QuAFtG5dscwiGO5uxkeMTuvxv/7QvgcDf8aDc9dWn37ZWUHVxIoB
D+aUJ+nbU5kcvl9gpOQ/gpvlUun/O2A7alt466LzdtghBkoLShLAj5tJoUw0jvZZWxNeHbPTeLY8
IkFOnJs8GXsItE5BSczo9lZy2dFxs0p/LLpCP3d7tZr+tD/czew+sVVJgY7o+NilNk8vhM9KQf/f
NNtHgxnCznKsFbqpoee5p+NNb4xsDeUFhnjJn6HpsNJkobEjXwAeL4czuQQ3u9/qEyLEcjeet3KD
/JqQ59HArv57hQexF3rgrSAJwBvc5y/9rebpiewZY8WgcWzK1fCxMpJL7VLYbM5pMd703qeg381g
luvhqBLx6PASn83elVCdLIY1WL69oCPLuccHmGvomf8S8Gy1tmc6iERiA8VGT52BFR2el+5q5Yhp
NnduORGgHK59E/zOTfjCUhRmvcR5ezPQ4Jmuz49JgtBbtNy2W6CcdCtO5iCPv8kb6IaNpTaQe2Ps
6rTGw/6Vg5Pog14vawAQxbjhlaWdNXF7+/U+NKFhiBW27945ReOo415HytQLurNQQD4pVaQ1ynuC
VmoZNiyAKaGS5J+GdP+11SuLCVenHqUHgBJIJIfeGAknIiMUsvskugb+iUo04iBPJJrFfCZsrImY
6XLShXh0GKnOoI+NvaCv7H4dc4uCeC8Hn/4KiIKo88AdWmRHUhJ88tHHosOG9d1HmbxJJLuSKCMX
D3OdzrcYcLQsr+AyjvtXht/6TYQc0LSmlqOYr1L/a/mSsClmqRlP8EWY1Tnx2Pf92q0Q2YxL5YIt
KZDoZmy0q0JkzKH5lSlQQmdWx4mhGofE3Htb6IKVIG0gG3ZtcaF0Xm03TIU4JswEPM11p9TX4/m7
6YtJIlwwtb7NPWgqfHd+WRNYOHmIL5moTq2bISb8KN6ivr/aJDP3/nDSvKUcQKdgchvuKzTjIlT0
cj1Ln03jUf7PMzl6H3LFDDWPkA6TOsN+LPQ9WBIt3A0IO+ejM39afQVniibC2DZrpoi2s6xdUz9b
e6jBH87dmKXmT0tXXm32BTwQ6wrmh5jEeM5bbr1WEBilxqdDJXhazC19y/rNJ0nNi27NhvYhLltR
t/g/J15c1czPnGMHHsT/y8b5nzQfMwt67b0JHZKaAsbp0h/vzpso+BDin8MUww6BaXmRtkv3N1rN
rxECKvFFjJrk8CFC5O0VaBydtMm5uft6bRkyqUBefW/lBVFe91iYwFa209VNVxctWLYAlUwszBME
FsdoGZ5NKAxptzt9psdU9VnJGstnW/AO+TVZkw3RD1dVFqwJV7yGo7bCMaZQmmPJDH8qhvs99pXG
6lLpN+6WtRmayPwebs7ACLAOlJTjq1e5gCZ4cYEFVxqgVCiNBemY6l53Pv0HJWLK5r1+bVwtSVBj
cYnpNrHMRU1TKCI8BJ7wpgal0hvgsani0qM3qcI4oeiMaz4A9tXOE0mIdf4BRcakPaCa0CbaROKB
Ci4UFjhSybR/gKAEiutIvEO2OBmhl7XzjPei0lhjyaZcthIzGVfyGEVCVc9FkGDrmKlqwx9h+gaI
1CULIxajVBtyCnlUBBiFatSi/WoauWNzPN+2S/fPrJsGsSOGE5jkEgWVBoUbWkcn49uc/pb1lwpR
BgvCTSoXk20UTQp3MD1loWNNbMdDOzS7hfDTo8dF9mA0i2lH3Mfai20tEoQeS+pdzu1ka8t0CfFN
JixIFd1FiwdJg1mfb3jutCNDfZvMqm75KuWASEDLF0upli2QtOqSvxD+eTDC22UCL0FxSN5/pxQF
ypDLKPQTwi00RhPPRd4a1YG+4I0ehCYJeUmEEqptH0JrbciRfJsZsq8NIJIRfSStnZsCKt7UWlfs
Fgj8YJJEPSB/w93t4+sODg6rxHk83bRZrDKjUZ8WYh98LR+jZ4QA/lVwW6g7aUIE5mSswhEBqDHm
RVxFZQHRFFY9Qqrt0qF1quKV2b0PzeB2v7MYzgrFMs7ubl4Zs/x6ZUsdlQYR1WKO6JY/6jkiP1QO
WsNpgM+MHy6Ai+hmrh+bTIJdKEpiSJwFv75tMSLRNCF8+rrBw8lmYlK8f7x38kn8YxT9EIPGSFq3
LT1jDEFpl34EelkVSWze4v0vnRtb61HShFZSZigI6YAjcOC7JHOp3zYUTK08GDZROQDKQq6OWn+o
+al0tg09yTJ5zj+sWVioXPWDU557ZrSYKO47mxc55DmzbxL0a1XRlC2ktvWOzhCtLAYN+9sFaOLS
r8wRIYfdGmIGc4kghzkM9Ui03hbC2p7Q74/X1LtFxJ7omsSabrNOY4fIvIMP58JzGTzzVMpHebYB
Z1wA0W3AGsGFGQUU3YayAi4kAD5yODa6lVJemDA+428WrNsBBdksrKvr94ldKADTmuUrWkeRU69l
gxa9osSHXoiGVCquNR6qqO1Bt8akB+X8gNvCjaq59Zn+2mX/qa1DUhwVgswudB4gQpMaTuCMzU8S
sygoL7XAgSMeT4i5rPXxjx4+vN97LUvC66F+OyenbeAEy0utFfRTcA2WCVD4OMsJCvlgGnsdn4EH
gDHSc20+zz/IfIAu7CVpT3lnAs76B5jXHcWCdh8YsMEBOTR5toiEPZg2xE4hhE07kKEXqqhvGYyG
2d6I+GQB/KsY1ZdTOc7NbSYnjPuXEoDouBWNLOLJGCxP1dCrH4kGeqgvHgfMIiy5Pvi2iW+kMnJ9
U6VLOyum8qvb5McLSM9NDRNEWLEmvRVDd4MtnXTZDcShglvgu5/xyi5t5UiZwuTrc8tp7Va+tT4X
tF2yD12MPEke8/C55kifW0e7MJN9GMfmt6whz5sD+/OALlwsnyrNe9302B3QuyCnIqQhBB+AogWG
3ULIVFG7kEWygKrHWOevWo/nSD/XetgocpklQCnxwcAkqGekn2RHwWuNpdiHyzJBnKhfv4dokLOI
XtWkDtoc5VWPRSxEQU4Chcq+mE88RNfLbKz+d5vwjh70r/Ojq1QD420HzUnPKK1J5+72njMimvzC
vJaqttNbHuANpQlASWFNtVzSiCZ8CLbeAFesu602UBmJ+l8nHt0YfCNsHCi5UGF91MNkozodFtpz
7CkdrEYYUqcKbAoW1Ur+Zt+5aIMRhaZrfFDRClPBHesy2c51wykjLE7qFaVRDbLmD3quhNIZtEgE
cDKdo0Sopj1YQq3Wt38k+KToMAxeicIUzFThgQaaFcX7v0gKnraLvLJC9AZ2q32G7s/VzaHRzR2O
dxmP3ADLwL4VZYLDEk3AbfxCmd2/8O3kXVesIAXFWo9qcGg3EF3wXT1xoFKzOo23PzF8Eqt2+SmS
qxg/yTftUqEMj/Hp2MxmSKEXETSR3bE+38APw8JO0Ae0bnfOStckBM7Yp/GSjjfU+qhv63oHL+vR
QBvOOGRxTs9HAhUjT6Mncm4+SyY009ZOz0X+yfJnZ95cWTUcuBrBm1aSFJom6rOi4ZZUl6hagq2Y
/4ZZZhmiAT1g4MOkvUGcLgVmkyfL7km456txTA27BnCpsQweYRgAG+vwcH5jHLrXil4WijNTgYDa
1zyrB13qLghoMQTWMFp7uvM18iJ8CK/XiKYIoMFQtt0Gs+6VWpA7uVo1GOw3Brb+n521lUUZ1ZLA
CEg4zENNqUBITo2bLcMIB56ecG9aKf6fqE9PZhUBno3VJ8YzDXCzzVZONJ17WU3xDqwZ1WjlLHh2
rm3icVOcHYv3pph3tB5TEuZF/7AWdxRjk5Yx4dPV4nmFI7f3SRL1XexT4CffqNBzs0SPKa1jxCgX
I71rRs1mjw3nK9AIsM4GN9Eo/ai3anUey43S/jaUU8UuA9vBv1qXVEzIyAha5gS98D2D8Izrsz49
fO1MesNWb4T4JrGEmbm5RASNwQXhSQHnUopPelBHQiPTRRaY544z4wQBAj6fk+1tfuuCErWEE2Ec
Fc9YM2XlAeSfd8akFiDIOD0vMTpb8WuDZR+vTxn2i4q0ZZCkLbirAZsWHRqcDrRa+ZpdrCGGQl3M
O7G6Zqhdih8B4LeN08xvjU6HMMSLrDFUH0vu4wCk51tUlP7XbWcxfHux9XSnsPA86/HlvPU46KKz
dQgEyd0GsoM7aF/Sj1I4kfIyZ25v/4CnXpwh3DIPl0BWIz1YB1w2GuUxMxMcLzl2TNX3NVo1R669
MiPXjbzdEr+Y4V8rxD050TegiNZRTq5uokaPIC9kic9wzSoGVQFFgOSKLFEy8nSJlO8Y2ii0DHvy
iryCpbJlboxsAWdYvrRHH1OTN82Zt8WW1YDb3l74t/tT52Un/2df6i6M0xL91t/AzVscQhbQmTNP
xIybje2d4XsAJ6BEA7lGBcOtiUnEYb/heCEEcIyoV7Kg3VuOBCd8G626T0+TgdUB3g81StlsmZZ3
L2KY2XPzYXRpX68TepurBi6xo1lczCbuWah7XLJZFakDq2YJeWuMtLIqwhXV8/q9jNrP3Km3PyUn
8XICW0i1ukH05o84le5X1GQgdZg2HmNJluQ2aGa+4r3PDlyIDXMowrsd7sSsJjzzIHHvFmxGJz5V
Usg61o44O8qcpktL715K5OYZiaonWy7dpYLViBJK1MWXYsyYMHRs9ZsXjc3OR2volwZi/jO3lfOS
FEbzAcnyjz/x7f2jopGWsEMH+Y5tizWiFEaeBZM1pOdYmPaT9tVZLoSmHYMqbtQyUhZ57vvVfoVa
+bduWi2zZ8g3OJIDHuIh8ErRcrKuTBscVAC3rZ846p16jONr/36hoIQPOyqougxCTsBVoBv69lx0
mJEId/9O7PUSRAPLUY/FS58hGqb++jo7fWOvhHaxLzCBSPzoTUj7pmTv1KhVux+e/y4vsIqTDt4/
xHN5bxabot6d3uCYR+n9v4BsuQXAMBbxbmFDbzvsQLiRHBdySH/QjIP+YrdkG99WoRwzEY/VTbt6
uJPcVL6EH7pQbpOaRBgV4kHfMT73LKFSP6bBZw37kH5UEIc9j1h7B0NVxZgWRxjbIXjq1rOVF7KV
nvupEe5AC4eISUtgtOfsUTzxtNJECCTBvXNhxhL210qXsP93pSn8RdiOg6j7FCNv6OC4Mc10KyF8
5bH7/arf3Ni5iCj3rb868pDicDyXyr89/lFU/hW+NAdAubwXeRJwo07Whu3b5wqoKKOTF/He+ipz
/RaZngB8lvEiW8eai+8fp/tqsJxeWQW6M9gdA/l2KMjD2EjkluRbU2ctEy2nQtmUvG0u2s1psh/U
cjXC6fd4gfuMeNxHJnLsarII7wkq68QTQS54vsdon0hW+Sg+nyFet1YHKnvsJL662oxAfoSw9/rz
PB+r93AyypoPnOTXIyFuPtJZ7yObFsw0pZfq0S7VdEe6atYefHD85MMZK4ljC2IQZXohUH0DQQrE
sZR6/gEU46NazydncpLilTzuS663yE0YhzNwnpxjKfelDVwqnOPbvVX+sjTSgWiO0J4eiF6VzFoZ
VIurpMTxp2CXgjaNmcsWAGOhUB4XmT/wKjELVUNB/i092BxyCQ3JBOZJmO44GDdYo5U4y6AYoTnF
shxMS27ce2BOQ+e/GoX9rTVf0VVTrFmxOXEOBm+RD6FhMmCUUXp3KTvChrESiS4V41UqmlFiFwI/
//lRltTxkb/uo9HDAS3PolPgxyKr/VZ4nSd1JZ7d4yIKaABZ8RFYvYT8ZVrpSgM9FAAZnqO1QvLM
RcX03AHTcZGfS7WBEIzqfm+ZodxTr8kQnXtQUDhLJoelf5MaiNg5mGDseWPPGFDsoSlbQxA8Xa30
f0bAIHCQh9R1/6X6BA7At6nhDhxiK0zZgZSlQHqLkRs9j9k3rbVXDvrYfmWECmrOPamALbQmiwzI
EltDHZSwuCY4SDgBUgl0coIGI+Va116LaR2SqKGX6lbWpAXILADR9PSE+A3gQVe1vSImz4gWuYya
ubwyoWmFIFLDN1fZpytR2I5vTHLvSl7QL6KkkEbkVx3+6Sd+14tKw7GyWLCp6PVYbKAP/UVYMPWH
m5uFrJEwvAkvIGghG+1EdKhjK1FjhG0EITZ9cB9fgwR6lo4MHETpYoxRilp3IuCPWHkqHVxWS/8r
+INgFA71vYUCU7e0ZWflE66XhqpbEPlfc6vTGyust5N/f9zidB4MpaDXBf5Eo8gp3uZUEo5FAWP4
wOKvWrstsbUwuyooWpkf55XQEg814/7DyC6wntdmb5BHQZnIf4hvjEi/pxseZ9TYoG2+mDJ38mOo
8JqPhIYSLO24pSod0g8t4h0dbAEk0DSJs2/BRwC6JDyNW/42WJanYtjwENpnwmLs49v0lc4uW5dx
RAGiSaYxbbdEIZNbRBghbbhUnOTAuCcGiFZBnVt+Dq2ES82LOokPS051v2f+0GQ/u7KPa7lTJqQN
dFhqVbjUFuQfLRwyniegJC88DWfJmmr16CnC24WRw55i8GEpXmbfu/J0zytIBqrfn1Ee5FfRkwfr
lJOCqJ7BEbtg80vTS5w78mmjwaqUgPO5t5U4+GKwI2y3rr/5WX/299tt3sUNEjZP7RnpH4oO6I/I
RTs+4/g4aZZXeoKJlW3TSk32zgM2KsjndHyb8SJC0KLAKfbxfwD3UfpiSVUJOpyqSkbPH7CCbahu
09BObWqrc0OJGcyqY6qwbWooxY5dmAkDg+ZSgxKJnsPwLcsyD07e4n6VywZINdNBFQJOuQZW/ENd
TbkZ/Sfk604mfOTCUo7evVtWb0Mt2WjxraLEWWTEkecLcM3YUqK4MMKkNomac7khyexsbokEYHMY
s+We4bbccT+Pzcjw+OWMcgBvprraevYwsz5DgDVhZ0+3YaZNO+XIP7b0x94+5gIBMeIR6Mfhu75Y
fe3kBVlT8g3ahTlcLaCJXCfEziyZI99lI5qUVLA8YSXx4VmlWrl+WoceUGXE4OzwLPvnNOLvn+CV
H0z5e/O9rwxDPZQV0qc1BYk+zZexI5IaErCdyqtqU0N00SJloR8BC5Eqgh43N3/SY5qlpSrdLEQ3
8GFER/kZ0d21gZLEWtm0gvm6KxgdUNKE63wYVxbbkRXFzDpAipa15oOQzZbbCj1Mzuhf/48FkNZe
VY0QOzhZR4otjf+7HhaAwB39rDRjkfxKtETL5T4CHStGNg1Dv7nszr9TLHx7ZF3xYK2fBqb/adTL
zxc2rpMxZKB6ZOk6k1/c0hkRk/86vlemJlGPZMbpiXgV8odkkJV1e21i0+79+51GXcRaJ9ERSFBb
oM+gIFZ/y9Q1vS4wEtd2gd5JZ4CR7mxgB7bpkzBDLM+PmZRK7nJVXCoSUGGiWldXUVgISR+r9st7
VjLXz4/5pIFUoAcjjvV1rm/LxtxiBV/wHzw5RoEKMWVzHoeN9fjeyFXBZr2utBuy8qkN0ydK3XzF
z+T8HXvjLtRjxlGNR4ZYMgx/ziVl48ojFgr74hEJ3Ua7JGqeUKZneV3q3j0EdRSrpsfl7JlI/dRy
c1qARkFITiMba29Z0xcP01LJUk4jsbOZXMXJdRIYfZoI5O3iuvCXCmRNe3vnIbJ0UFol3088BVQM
CSCfNkOsr0JiA/g3VszTr4O0zi7RPxr6piIRkeyb4kUFOr8xBqz+KCYulioMsfoUYeBHW29j4xwV
jpa7RvJ5IoxQXGFlqvFepSwQHqUJrYLlR04OkgipUVPrlqNqNKhoF96JRySVuramkaO8k6FVnIXA
sYqqnbAt7rYsO1urTJfCOLSNB5PUR7WLMYSbtUD9CmExzCbG0tSxzi/AZV47tF68+QJSFPFH6L52
KY8hhe89jqgEci6xL9vY0uihtxTXWdx+q9RZLhaFSZnBZgiPdP9jSHoesVVgQw9KhDSPNxl/6LMR
DHiXpAxm8jxgnCffqh4I5UjPQCOwRpjzmOGKJH1Usbk2cj3tFyzEocRk0LRyYPRcwp0vttyjmtxk
jerHS/yQIfMN31xCmVOS8N2JLzFfka4ol2rUIRm4WMt+9mAPhKeH1f6T8IFn1sQK3fqwiPlSoFjQ
AVKYP3twGZsNA9hpZhFiTlE3VTOfWtCjXkcy2OwysiFa9MsNAlHJQnXgyWxwSmfJct0XtbEsaGOD
o0FhdyzzS9/0E7d6efvGWK9MAQlKcOEiYQCBRpNQkPbwwJ8PagKGa8vFwQKpridKYSogxvNb2YSG
g8eUw0ZirFV6rCndtBHqkvRsfV3Xdu42XOijyXp+h2x+Cg3CvcAZbkIJBgc4yQVpnVaKncy+b/id
gTs0aJb4YK5p/DkHlgxcyIDNnLRgy5OJ7LTJkEt9m18SN5lXdot529Mpi72ZFwzYqJ33BxuUPRzA
EuqSGDj5MPAT3mk6MhHtS3WydeVaSCzW01o3jEQhsXLeiaKMe32VGXCF0n8VdHRoz2BLKsSz6pba
4UuwEYmipu03SxRrRxTtk/0qEnC3eP57rcVGWL9R0n7PfPp9hl1uNOl1JDOuYIoDGfFWM7zasX+2
tpQFOZTJ5JHJlNyldpCK9C6MJrqKYJKU8ox327yGJgVUKw+w5ac/54mTogz12pxAnyiUnbfFkIUD
w4yLgcQz8wF+3jNHFPt/1kB6BZtTZOdyjHfTg68+nqeE25DK5RA76BB+7+/pwvADZLSH68cw2Gwx
mcCxpQqdUm0+lfs9OkfGB+SLQqR4s2dIkzGHp+DDQBARm0fbNjejIRkHeWOh5IqBiazabQdVheHw
fOKJDIBOQbBKE3swdahEiOToku5bT8KCn5cxdBlL6Xmz09P1WJF+c/tBPcDHY3SLgCcDGP5M/8Tf
Odmb+DqpdERdZSIdhnM/KWYhAiTJ1q+6zPoFWJZCLuNTvzBSeb02EFEekZGD7+2U2B2nTMS+LgDP
1iRlZg52qbrTgnm2NG6FZW4M8MnPPOpEfIu7x6a6fYyPkZMKD6jJLFEdkS6Ln1Uo7KRRA5/13jOp
ztcIneBh2z9hkkgDN93OnUSK44PvhykqmIKI3SEODqu6NzReNUOpH+U40phsUk8Iv+xhrqzgsyUM
MyJ90Br5oyXjdRmeO8byjx0YLayTxl4yDupcMF3B8Vn+bDP5yKC8Kuqkt9VN60sJq+81hMBYJGc9
1wYsHmcyLvj1RLYNapZhn1T3XzDAjGy3py08ewSDbM2qfxec46d/3fRVG0Fp4Pj4/3RqA60qt43c
uCH6DEppGF4hd5lHeewCR4tqPfcQBKomx0Pd0ZKekDfFA7oe70grIQNSu4GXN4HVnWDq0NPZCABD
HIqRYMKB8AE5GFwBu2N+/4U910d/qOCyqY0Z17FBoIsecSsiDHN3iBkfkr++/+dghNWNHgVAcELk
3hpZM2XLbY+PGm7wGJQvHNCFICv1lGSKtjv1gps9n1HXs0Bu9jaFo8rjca9aCO0O2n/2LrBWTYOs
EaQfHGWHSc406aarlN1hPTENGCbAsrT15rfk4ydUjApj6rjjRH6+8qu6Y/HYB6W0o40wNkVud/K1
rzDhChz92e/r3l60h+2ccvwInEcTdim47WKiWcQ9XTmoXOf3DnH5dJJmdsBluEyBgaJ1gzuJU2wA
dA3EvbI0CiSKuuB/hkHyJM5YMcs/Z7yvuU+3pdf67urPxaJO5x4t9OpLLK73k9uEO2XOJnhsQdii
qTpmhFnW3ErXFIYNcnwp1tyb8EY/zDddwHtUHP6Esi3bNVjAuencOUoQn231rlpWz+djEMFuIGiV
v/fCFwvILF1N3/tQFIi+ljamsPXZT+/9/rCYpqX7sLpieusV3Ts4prFtqYYwRo9ze2D2N5LEoSY/
IIN/BUi/crxnUj291WA6mC0hISJZqLAo/i1qxlHXN6KRwf293ohyfhzQY22wMIjEQNJ3JICpqSW3
4kwOvHssgUHR3PARlZQn4o/acWXw1qE/g5o5Rv9sILkOX1In3lfcwjkR+wJqxOTjMrq0eFs5+UNT
L/5qtBr2tWWPgoRRoYeUvlKStzi3ZR1RjGSvp06VBEbxjFuH71ZBf8h4VUVt1azw5durk3Xga7Wq
bNnZWw7NkIZs65glgfWlRkcsj60nw0XwJs3I5F+Zoe1fllzPHiTKonNkCEOaKVGT3qdrYCu03crA
2j0AqU5jHNqrIe7Uk9JCACZqwOkq7AwUsNvE2OexFH1vtr77ndqlpv7fuytihIVaImKdFLJwCfZr
MI04gJxRRHEUeeK43Sb4wIUKONevo3Fbqus6G95q0aI8Aq8SFeTKdTLlYiCU85pw7qpi7LveNba5
oRHoRylKP1+tunzlgzWKGtioWLt8QtmqPiWFwKFforYhQzBL4jraVIYIEOYRHKPy001s3LyrAgS0
AWstTORu4f86BQnr6upsmR1S/tkEb8dGmZIOkqCoKXECn0g+fmCUDgOUJb44RHII1zNhPlZLjK+I
SmfGAIwFqULlPspgr5wbsI8dvpj4JnHN63KHDO8I42zkLMJ2zbiB0QiSrARoFEl+RT8F+nKcUfQy
/oNhisw0tOM9iw9Qh/wBUWyhKq3JIw4eWv5BnVyg0uQMxFqkqau2E9a7xaPt3EYoD+407I6A0KrB
j+x6VE+q3dQE9Gz12ckQIaeAZdNbrb76oCQmddIw2Lkaml0JkN3psBMAInZ0t+V4dcjwf+O4jnF7
nTTGtQfuLCpp4baNtcdTV5dmnflMBRnT3o7IPings1uT56ppveOWwOtgkQHJoRR0MSL8BABVizaX
1Mf7785+jTDic0JQDCUh/OcowFkkHv+auInqAOnkrVnH0MbonPCfn+3/qD4egk3q66ki9RW+sxB1
idRjNlUreWyfrvHF1eU87Da2NV5uzOfUK7W5QdpvKjMPQ0+0I8c5bmRH0ScrgYHQcmWYt9sRYOPd
BZs6rUq3JmYNlKUt3O0NQCElH/h++K2FxoZiuNxPhBFeETrIA7UKzuE2cJjcQiftx1dh623o/gqF
GCi5FJm2zQwL4SnaK2nnJ5P2XyCoStvuejeMcs13DaA5W839q+eSVLb+udJoVxNuG8HVrM8WIJzd
/r9WHfdo8iM2rt/ikMkUAzBMK1Oq8lweMQZTr/dTD/WlPEcPTc38hgXfqgjId08AXziUF1yYK1kV
IuZ2fCrlLE0Fr407HPRQJgNcOyTW90/e8ZBNlfm2oFqgdNzQ8Pmb/5KUc4dmAslryrcGilBoug5e
v7ghvhuiAmj0mU7bWboMsbJ9OilIXvrG4EkBh0H40w+GjpaLk9Q0luNKXcvBCIU7A1gRIJKOkPOa
BzitwZutuBVsnaBkan8nZ+dXA5HOKkCjHNOBxbVy79qLJHXVMX/ucLNGxK+P+mMM3iXBTGt6QUnd
by0mwNdcqf8kJOfXHg9qxG20C+vpxEg3T0xMzPKe5pN6BOyyXIHkVPB+TVkhNeKVEtolV3riaAqJ
f+CDxOEYyEX6YpDQ5d9BjnbjToOD1fdYCgOVcz1qj2s787iy+8Tgoimfk2cBLa0u5aYvmBJWe61Z
GxseAhA4UdVDqGgweLiXsGuCLRPVaqz/ei/P3nua2+MnMoh/9HINDpY5rnBoRB4X6Szi8xhISFsR
FCwQrKCLechtMc0oUUS7/OT90+eYTn0TbCHXC2PHy8BOJQRhfed1Yy5hhudxx868Io/LliS7GMDK
N1NQm26R+LfJ5EymhwV/TChAc9lmrwgcXuqY/6SZ+yONEpJ0DjS4Smrv6yFVtjRA/VxjCCtZRn+l
HfNNZbFSMkE7bg11sqxapJnkLYC8ssztBVWkgUj2N/P/5ngg9r8AiEdUWfZ/Au0Eli1fnDal3A/s
fSgsFHiHX58SShN012sy5frFASWbD/xmVE8rk0NgMtuVLAUPSnB1NRK1aeKoWBR++v5kHlvPaZg1
yV1tJlizSM8G6GuOB8u78dxTiF3gDJn8Py6HF6o4wQ6bCcx52l3FdxkKjQVGphm2S24+/j2zEHee
E+uZWeJIXxawxBx2kVe9m/DNCQYbbP5/BxoZE1eDuQN3S2m+tkDEYjYnt0Pv5U/5uCVUmkMLUtGk
cRiyynkbWc28JcgJLNMtuf9EwOu9sm8TLtJD+JQDTk+zzj9TeW9BpOCSdnnXOCjuACtThZ9YIEnv
OI7RHSBDyebG5LYchcJy4tuJgB8LjRefN1uqOnIavN/01u4Lk6Y3RoApeoxLzzvuwMyAVeha9AWV
L5PW9z1gK0Ra3D3R0EKJ8YR8UYRqba11Pm6HLsLAOR03jvU2p/T3cn6kgc+krIKkR3G5UZHYjAku
W7U3LyCFQ14FhTNDRkwhDoLeofA2GkALwx64ORpw78aqV8gjCPFMgXtcHIF6p1wBHgw43nbsFkdZ
MeLKOE8lhuBnTG+k8QDR/LP2lVf7gsuy2ddvYMZUEb3nHS43oiS2WZDa7R0Vr8wOkzM9u4LUq9Wm
O3v9dJ3l8h7hMsC6JzudFBXkPD+4/gFcTNyH9NJ4Lbgnh3HmWOBQ7iEhG5r6UU3FtyiZA4eLkmK1
Q1Vdw2We9LMCxfgQyPfKyT58ucimoIZg8kuy1mT3hxuuzEzt10qouJs/DEtF3CR6vBfjGv9BHKNy
V64mA9EWYN0fLTObIW2l2g+dza4MU+gNNkK11PMNI7RcJhIe5HOofzHFcnKVJsBFDXWQtCXaLCU/
KRPuotsdyahAOo5/MxH5UVStMxvn3+8RekfnO3F6ElQkN2upv2b2nLTBqKEhfnGU3Oa8OMgRjsmX
TRvRrZ3Kuf+rrsNCg8wlTr3Bkd5HOAKAVOTA4q64POKil/PCVFGcFffia45VB5wCEKq7mAB5HMDK
/kQB5vajTOkvkDydPBkHOsq9Ekb+/qsy81/j20HMjraqpFkBnXk3EuCXqbGnRAmCioFaOe5Fzle2
qMBrn9+JasWcJSnt+zB39r6qV0ZLzC3M+RoRDQZgHHni9/AmuALWbY8HFYvqTwfG+1ZCxMvReEcF
pUpo6n36EEq14xnGqSSCZI6wsguoY0XtQFSXMb1Krpq08tIh9RQLK9/tTJxM7ro87PDR4pchmlTv
tbnx0IuUINLkt5RY9m4Sh6E4Ig3iZn24AvjuRzF3dyZKFhdQgtArLPhQo3RHThMsmtEMsUMFJwjv
Ap/xL6mick41rHnsySvrBAEGlmMNkyRC4oAMDX79ZnTHdIgmvR/4RgGNWYBFfZvJrYORRvjNuNie
dhzw+fnYEpvxsruulfChGkYAu2wcAa+eRJHzNxbKG3IgDDT2prDXZccYAFgJF3xg6JM52SDioFvf
VH4CxlRQfhAFXxK9AYPeWAlrqsAuGlQLK6AnJ+QluBo/P/VUlHL+Dyk+i4EMz88KVH0eyktQQYTS
/jYH3e7LXhuevT4/uhFjT3JhwnCTOV3PiCKPdgQGSVLy/IEVEiJxQLM3Xbv1YjQEvRuhuIVxmH03
scLFhFcBmnDAEn/q6i/2JNGcjgA5b/zwslWdCdnM8BZk7dRice8DlUUtmuRplNobYWQlXPk0kQ6S
UKvx9f2hWzu2vfYLKvoSo/D5zPEGCcCwIlctAl6pdqvYBfvjrzAKrvT/ODrMwxpcVUet93b2XMsf
nZ/fJWig4XEYBJCe8eXgw4xmV7SiVka9d4RjCe9ou3ZpZyc9ABvgsfeR0JoJo71mnQr+P+raAedO
pGndrRfuR+1oQe8XGLZ3rE2vy4x1bn+/QtKAxaqltMP92YtuCe0inTt2kx77lyYnZgPnX/vDrbZM
i0zL204WlV3WP27zibbbwoPtpFMHgftJCUzHJnmx8IlTb9L/vH1Q3INN2zto52h+8saPGgTQYOQn
8hWHoIkus0enHx37urtMFYFd/jYki5v/mXkmX1NFO+x4FGxWRdTnkxdfrWziau69BERLHUh8m77s
GbAju+7U8yZ+b3XukU995AaVEYf7PPWy8lcIYVqiZyw9ayU8knv8VQNQmEGFYRgK15+g0fCZaeym
4qAOX0P1rqMlkoMqJk/hWgoX1dbq/wDxryAbbRllZ7uvj9LfyYDrwczVf7nWkvdoGLJFbJzqQCpd
KxdHkLix/DdhThurq8mg+ITTudqer83VkiEE0IxeW8gi24t7eRd1Pt9yu5czqYLPXRlnHhqVJii4
xIxqiJGCvx/tFzqVNJJD9qN4KiJYHGBJQNS0TwCp4DNgIbAEYhFHna0cYKmQX6dYMghWwuSf8SzN
3n1maAQ39ojUg7Y5opJAtrtfUqxJHWhWq28OEUpnpUUUKb6RM6Do0doYExJnf7+yB+1H3pbN6hdT
uD2HcamtloLiLj0Kw0SmnIbOoF0CFPPsOzfPPCmfrbavFKiZDG1U+IqZayCMenRm19Ac6whg8tNX
8L2YqRdLbchj1EWQi9XpRJJLezXtNM9i1kngLIrY/jybFn6ZeJkBwoXNYCqORaWDqg0ZvLnCuUAD
IJpa1gGov/DGk9DJ+IrC7L9NmMKNbhtPUS1wNgMbOHkFyOJMqnbXr5U0Mr0dnm8cftC6zpj/vsYZ
roOaY3LmxBtKX8NVBX/bJzvaXnNo+qr6EqE7SX+A77rPUZeGZO0naNZt5T9qmS5uY8MG87sZZhut
fHN7CZq6aKN+NynbPwYnGpOJPyXABbeqhWpR92SrkDOQjwUCxkncLbOL9ecn6JIN3G/eYGg3mqi5
CFJ+686D7Mwj+Amz6Z9Jzu/3l3bKbsd7xHrgJ4VuTL0JYBKm31V76qJbz3ctbhQq+ekz8tq1Jy3T
ES6z+JRJpmuhP50n2dSpOcfJPTWvjas0MQU/ip3ZrxYpLYBr2jz5BoPgbSLTDhiDXHgcp9d1I1R6
+YJQtiHT1MzwMmhqe3h2g2kxneilXbVk0SxlWTtdRSp3uoWr44DiF7o5tPoPhG+XDk8IvJK0jca7
zq7Lz7CPkwNEkxEeciJF6xMWrjXmSmxU20sPGB5yHyG96fPOE6R+8RJs+Qhkyi+sORJt3hiow6Og
V6c8KdXDe5eSaYDjKLFgzMvjFM7YGLxyspoqBcI+Q+rTd1xHliAWm4/8t7mLei/ki9CknD362pl+
+zxxsONq3Dy/hQ4iqXKwYf+YnkIxX2tlPaQOKzfth/BIHjeVZWpHT8XT2DQg82M5UnCHbBaabdiQ
lDBoXKct6/DNF4QI3edhGEqbW8Kghoh2EsvrY+xL6KJXZD9tiHcvWlWRB+Ke1Mszmefh3xsbcRU+
RnmMnQZgkY5ez6MlWvEFbrn/eEXhtcq24HFhhaO9xMsyPGR119mllSYRQszW4hQ9ZkJAtu/PG88q
f8HqmtLYFXQBm2IfEiZwdn3u7a3Qb+CLo8r8FcCj/sOhCnVD+g0gI4Bzqf0U3IG87Y6QC+MmzIAb
vdjJgmFLWc9b1yVqfoMm3fsLyQmEeO3Vto1mjXjlBpPNpP8RaB0pT4Rns1/7KzjLbViOtrqbbJS5
eCSnGe27kld5xpHHr/cWedLSt0ltIU9OWN7Pwe611P6E9RyQlRZPAh6vahquAFvCWZLmodSJ8H1V
j6QLwbLwp7bb4vnYMNsbprZr3kcFnL0hjifuCVq/nxHh/0M6vQni01eTOBKII3F6oiRVRQnxcHpG
3rMNum9EwO9CbQOS6BhEr2O2+1YFArmp31GSs6HxUbjFfbTblJgIqe4DrY96R2JZTaeKLNBvIBhj
58YQAxm6Y3GLQCBg26rcl1OAqWBTQuPRtlcs5y5Amjho/6PkBg4yXj1DzLf8r/jtRYED/YdReFyM
3fhoW+3W3MszVL7j4t/HH9c4UvOQImj70X6DOK8YQqNE+CDxr0dtAGmO3ORY66PG430dILtQb1Dr
mShtwpjpWdYwBqL4hhFW/MrSZLLzjhFocCLIXZuhEwhRPhvNZljhl+faGVUgrJlkaTAq0buF55Sv
C+ePnteer078l/GN5yzNndObHZPUKf+teD98iDOxekxvYnt+JyeuB5Cv/UfR5cnt+nN6PQqih/XU
HBJi/KoBlfPrwjZUSO8zcm35nuhLh4IO6QjfHRib2GU8CgWDZsABqIqEI8TyhHjjP7dK+T2mpXty
U3WHEto33vTrjTmgVm4d6EJSfumAoi5/d12p8wB6HEEqbuqUPhiNeDWdpiEYNX6QPoU/nGF7ybRi
udddReaqiLz47R2TW4WnH2EnlNqocBk5KgCzfBTuU4y3xZQh0CmxpB9+MRWWcvz/fGT6Ejtqx2LC
faMJsnQA0CYl26PoX0wdVp9QCH39vBEqEzGw9sJSaZBDzfGF6qnIcgRDxtwtvdZ1kLwq1K8fOw6c
smlbLBakgXY7wPKAGzjTrsjK/3QQyxEFbd66JUQMSWeNl7Y024z6w2ASK1/rcg3Y3Gq4N9iwrSg+
AiDoOMFI7SxfB4UeD/Dcow4ARlavF+WpG22BR8Y+B/J6jRwAEQ12HkEmUW1cWABa6QlKJ78t0LKi
Nq80PQlqNoW50DedXkdbzEtbdcuBmkIKt4t5jHEdNuOBEd8hMpfMyYYqHN99TJzvismIQ31ZRYfL
3+y213rzMR3yeRJYFKp5C1KQ6sn1dx7zyohEVNuyYaDNGvNWBEyQFKvtQoULz3X1547zqAazKYf/
B1jsX4OeSz7tFKVGwP61/aeyae3nL64gdrbErFx2GypEuKCzUH97XbDzTsD2HhWit12pwztoW/A4
2v6Gqg0ldwD69D7rgdpkTSIvFmSBML931YY0slDWq2m3Nr9co579/Yf7cQiI6af2x3VlWetgqL6L
mcNd8LXbD8HZtSGEAZq/ms1fLrpapk1ZSjyZAM4wxwYu2X7LHfwhjIBeDxMn4FjY6zhYJzsaKHez
vALBJ+6me1lCE0K5lk1JzU8kK13sMn/EaJ2MuugzLAjLpi0b1+I20EpOuwh08Zrl2NVGLdyzb2Aw
xgPMKSOhdzVTDqozeoBarb0bui+Sx+AxMwbPtmSBl2xDfmy3xugAXHs5qmDdLmm9v7LXac4Sv0kT
uwU6JSEPB7x4lwvTQiIKnLKyxKoyN6unrT3yCefp65yU+F+lGV2N+D34dOJPPjt8SZr07mVOegiR
vH2BdsJBoWmZySA+3EabmeRbKgTFqWtCOiNHvZq5uSSjA3PXCRq76c+UubWWn0CxzoTWXSlrfB5Y
p3d33NWQtGloXr09Kg2QgPr+n/aUq2Aa77h1iBzoaomhPooU3jWYmyZjjJI4KskR/ABZy/zqDrR8
I7OLofHW6V+edaKp9cGi5wvllyL0a55BlSQvpz7zZZoBQBs5fWdsdtgrSAYxBR3ikMfrQHntoeLG
SYlntmIsC4uaQd19xpRM2CnSTYVVZRtuL1ahSS4/AOIUjj+bzuV70ruklvHr7PExlZrmf+THQKea
E7MtaNohJME9aFmwHjs2ikPopzN3KpaSd5zlI75o9VedUSG0/a7kKPbm91AWDSWFabqRDtxzQ/WX
hD6VeZ4MfBM2Wiu2bDDy7IEqOA6BbYM34Rixdd2rd5P7k2odtSw07DVncVei0VLdQPTcLTdRkI7Y
E3bWcMY6u3g9stXgVkjm+Eei76Vk60Q6qTLhULC10+ERamstDD3E9UeX3yJ1vj3JL3eRgEq5LG7L
qWFR9rMUstlqHuErkVgUZ7gyM0UIwsw2Hk2aS6sjehSxoMi/ObFmYv6Wf24GJjCicRmC88FEhpQ/
CLcr8dtkFOBfpa6cg1NZMngYoa5mc9UFH8ExoUVN++mt4L4YqDNmqy2G5ZKLCgVdINla5os3geYY
Apjf/mHcs6u5+Ml7z8aregpIMMcEDBp78mEhZzbTA6TOq3bJZr7ZFPk7CTR0cd8oBZ/x8yMHNNzX
I8SpC7VO6v4iVc7ei9nIljtKJ+hOndzYkPrcTc0HdBnT6EYOHQ0eD/YaoXKBI7Pt8VTrAPJm6gO4
v4Fl6IJIhrzz4oMRr43ZIPfb3W2eIykz8HGVrQxTn6iAy98xhTzzsOp+VBmKr1ksB4lpvVJoPxog
x0fObCdj9F0wNtzP+MLNGMJ//RkXY5amfenxWmAhlUIxahh44kGFb3hw6RKKyArcJuGD4GxyJv8N
KcgZc3eA26x3g0qp86Mu8QpLCql46Folai8oOVuzo1gWaAg64YjS6xoBKh+nK0SUmnBFvSA8t0Yb
NkMp12xKh1F09XIJ5M5/sslVxs6sgv0yQgRQNrUOCQeASlGySeovDoPOy1BNGOq6mRAspUicr57a
28gPUsG/EcOVHoyH8mTTjL2Kttlrpt0AMIy5c6AoiGiGhazeWnXpFS976Pe8RflPDIod+cU52kQk
3wJpccuFjK0YWpXwPmyQHaxoQiK7Ie5Vx3r3/NzBFGh1NhWW/nyktKibTdT/LdZuenIREwXTXcz6
z+A01BIbZBgxTKgusUxqKElTCX0L+yPKQEolOa8yBgf181qamwpcdsyfxm19+gj68tWMAgBd9+WM
ojTBASjUDf+H99Yc03IjiFFMXdgyNwjZ7YUgTU4NNADSEsycB13hBl57m8ld5UxDbLiWZ+eMtgoU
nANCpNPY+euRVgTfyXowjz5ArfYPXCvomHnmloHNJTX2J0+o2fRXYpc+C4bP1EU8T5uK8xlaUTcs
FX6/Mjf1Hz76DFQ5fP0KOqJCLkMhxMwOxkFeSObbTWanfFsm4e2952EzMjoEVJU5LB4+AgguTnSQ
9IbXLLWaEEIDNHzrrIRcdnYP0ds1wJwCS6PR7PiOICO+9NN9AeXgTG1anuatLYbPzmLCNDuP7eoG
p3LB29jbIE5ecdFbLjpNpA1tBdOHNl650dzUC8iuNHCIHHJQFXEhZkbKe6q1Odb7cWpHntyAHIPj
dZQvGrhKBAH7MtsNM/gejxxKJ88/alBz/UWoIT9rIcClgDJyhUWQsSzu26lAGtXU7vLWDFeUf3ZV
j3gy78fFovj/+gSAJmU9VvGDVW7oJAj1jLliEofEp4D5H9DjpexKe+1YmsViqMg2d/oc36cvSLZz
LECagkCBS2fjY816J8Hje1ICqq+zmM/l0gACWKeUwx8US3VMr1qhJpN1y3RTEs3KNr0PndKF4CRu
sX6jC2CVXfy4DpL/B10m23iM79ZdS4rAaHgo2JaZFCyTRCTKuVAXMc/EqFvnUDaFr9uL1N27knV+
C9V/sRHjVpmrvBJJs1b+/+8bdp7AFmFOk7Q+3qi7vmpI+JrvourxNX5Wg7LR/iLZWw8apWYHEii7
YI3FwNJXOUQBgCZZps9AmdPbOZEZv3y4AXDVyo2fGqJ8wG5fNU7GgG0g+gVj4cY8rdqNDuj7Qe6I
LcrSnuYwnNadMVHsQwVeypH5FLWzYnsZ2SWbBdxU+5zdUvNwCzxWLce4RQOoDR+6xNFVVXQYl5Tq
niWFUEWm7OpPy/uP7gOoFrbVSio12LSV7lJAqUAZNRQ79iG9SU2UEfbx9ex0iKXXi/LFyjHqhDAB
9u4EaKhzR1df4cEKTyyindo2wBUP6X49pQgvybKxcmTmCzIgaWhY+yKeZh0w0w/n0V2PdUKhEDd9
5yHqciZyR6cphK2YBC/+yLUT+MfqWiXchaAroB76Dz3v+dE4M59B4CXYErm05pd5yEhF+4SnSw4C
pEj+95YD3/OFhG5PA5rDILM/pDyqn9uXckskg3MkjZAAbtuDq5gvf+dkvcZKyi8BakiR+RBOALbq
Jvzh+IJYx0Capi0kqKFx4o6hD8QvELB6bcbzW7Y7cmChxz810NFtsQV/VYXd41heKdUH3JlHIQ/k
8fSlJ6GPIpEPtUN3B6hhd9RdUocCaqbHDurtc1WoYJGgy8A6ErpCojF23Vx0gDHQqBac0nRgXfyD
iEHlrLXEksXOF4SORalclq7afMMzKYFMqJRHEXLToyz9nGJuf7EGh2nB6qBlB8TD9fbazDuKuzE3
2vSd+OthFldB2ciM6ZKXqCqUVTJz8PICu+mvNaK+L4+AbMalkig6JunuQ0AR5nLSWZDeteoMVdYs
5HFv8TgDJqGkn9y5nvNBr6Foj47y1QFvT/4K6wV84y1Dw8JMbQ7XurQK0/EAvslTW3BBxc5+Do9p
lxikXOw4oqzQnCBJCscE2GyiVsxxpUloqKcvs5+EujER9vZjtvZGzj9bOcRS2tMfYEhlo/XJ2fFi
fXHe1GXc3vzelEQaceAWoRlJKbormwoDJtUCd+yVZYhg6ceYttjWmbqxv447pOWzlzwqrLYVSVJp
Adc3AlTtMg4HAxw4qaycoFIq4+xsPtezNLgkHNU5zIU/rneAd8KuCS900Yu0DpqLugwGVtWONk3f
FZnAn4TNqcfTmkKycmE1amuS9lC/6cjjtWYLPXgP9i4w8wpIPEJZBHMHl65rZ3fHZTGSD7cdDzu+
PFUtEvFcZE2YyLB1olboacoH1PXE3uMuGcl3wjSatTQFev8MsIbzoDeDKKyHuEoRFIqpfvPq3Fva
rsSA0tgjLmgF2o341ypJdvoUtKGgiOObynW4gpNXkwSyDLlks9HkvDFfmdb5JZ3GRcBwHQKglhnv
A6sWm/IHYEfI56huVtKwCRZw7Qn3u+32kCnbI0OysFML4lCF8+lzjYi5mJrYXEto2ul0XlirWH/0
Y1qXe9cQlqqGz/zfm4BAp14eL1tD8EdWCqgMJCM9JBOGnR6HpXOuA/6LYy376ptX37Z4ZbWQHrMH
ZB/9De8jeuz6fhXGP3Jz12yUhcJ767999Jq0I8CL7A2PXiXyDckU5tFaVf3APBwM6ZFAs08hLGuE
dPpvh4SLHmxRfhNtWNFUy5OZ/o7SSorBZveUL76FZsL0bgRZ0Mj3W6tnMn6oOkG9jdXnQQmWwki3
xVBrH2eIHR51sjVp+ilsjvau5wR5iXiHAQWjm1l2+SvjDi8BNBGQWkF+3TtGHwMQKLKMy+mlDzE5
n2MRP72hn6vB350L0KY2aS2EQ2vCWfCcP4smQuvMATNOT12dbYEX157BLqq2BVCGKs6H6lTXGlSn
VaBpvOkvM9s9EENgIhG1McRpqwfWlL8u5S84DnFuzGhSwU4qJZ9zFXzjpIgBESdgEMg8/sBQKRVW
WFpWl4orXL6iUEy7VvanNBXaIC0IuPWAVejQZVQ4ZZ9TSfbnAsX10g6HXqFiR+gBOA23II5Y3/nY
Ugz8ovFTip/7bSYPkRX13KEYT70tEhNggsSSJ7eg7DXtw2o2bvd05aFuo/7BA8hTcb62MS1fYzlJ
+pQooTqs974L0/TVgHHd2lV6EPUh8gkEv6bjR0zXm4cMeYPNEBomoertJ6VpTD5Dz3qBXBvZqAbR
HXKE2VXqR9hv+pb/rsSjP3YTR2/QE6g7EtV5hVP3ZByWlKWjYtoBoWdYLUb2fIJGkpjkiJ40XBdd
ZsN0n6Fd3F18ujnP2fjnK0ebFoXirMddLQFx42gKUfKR2+d1kcHlBggL65BBMpgDNo4HC51ZE/s3
eSSyZr/OMfhXX7FqzINBzEbiGkTS1wmnSSc6wKohN32oFpO5VvsxVzkxR485CeOngnFXHZfCHnKE
h4EonX380Y48JSyO8e+YRfwoRxVN7UGaLVoTQROFV9/ITgXyWQ6m7iAuUG7Pc3vTJPwArlA6IWyL
38aIZNJeiJSaFqIFk3apmKYr+75glmaFINb2Oq6FVXzLLB5ksOdatpW6AmBSFpapsv/cr2mmJRIi
DHb7beyGSywq9D4Hnh7HaHG0ymvU9uWyDZJHj0WuWmskTbhsVtWSXWB2GJj/RCwHSRcJkUsGbHPw
nhmu9p2K6P96qJuM5o3piQTpRlLZdNW9zuq2vjjO3sLWVvNBsWCYUEJ2lHqp3Vex3qT1AUqVVxLs
VdCn3awqA2ISUwjOEndhhFAiIqqSds/zY8HErcwndar1fgN2wELD3fJyqsNaKJkNJ+16irU7n/7C
tgN3qsLcrTIlu8y7mJr/cmZ7K0Ho6UbSeR+J81rNWSAURU8lEObJBKfo+x9NXtOfzlsnfGcsNhnU
AnPG65jXKOLyPilDSrIxRY5xh1LwG42bPiQABbszopNZxEU3ABKlreHD4xJ655YCP5/uBprsNRAz
DqDvG/niTtTTOYArolwNMIzUAfxzA6MJvI1WyrvckjNmacglmBS4KgYxkNlANuuy48AOn20Jepi3
oTK0adEt8l4d4GaMP4zM1cKQITnutqkRTZhu320yqpZu7inz4tyK+NhHKi5SgBJ/csqSEkKDSqMA
WY28q4WEwwHUjJxGJacSJclKjGyTBC8OijKBq9G6+rGTtn+yHqMDyOCgSQpsjtE5eoCc8RYR1s1D
yCVPJngAXuUal5cwwUyJj6oee7j4v5pbsIUFt+/b3gFLPLaz0Iva+XbldgrxduWO6p73cIiCufq0
foHZfWe/2ZZnaQ5RGQNbs2t72RnpUhNJc7qme495otfzipKHunmiZzYm+0eoixCNGYmxhnEaTUub
inYnqk1k1lyUKKQsNSbqsts3EpWGAy3j+IX6/D3KX8Qfuf5JeHe/1ihVxT+nne27AGgER530B3w2
73QdDXK5+EU9MPdjHy42UITQQ0ty7lmnqH5vePUyNliLWl7oV2UPi3abwwBH2Kk2RFSfT+9WlQt0
G9MJ0XGZpPTvDAMITY2b0LMFQsXAoyK1JivH7xfs6wFMlt7OWLvQ+60C8FB7GZUNipWfL1/yY5zA
gWUCv3u2wnYD26vbWBGyIpQl6kKoRRMzGdKVlNipIhYnKMDaT3Kbr4TzEn95rKxmTCkLX002D6Zh
kEd1+XgCYs3DdODWfqGNKJdXS7yIPwq7wyIyPCs8SmZXe44VssCi8zKq1KMu7+yZrMCjIhZVEmU0
XE5rJIOR0sIzWwXViSR0ObgYbPfbFWupn+TYAh88gROTD/1QBaJiP2cNv87UJ/DkEPKFFnaAT6/g
vGtQDurag2bP2mAlW9hwJWXFlButnShxwh4ULUJ1lqCdt7teXvggCWzjcKP8O1Sa3hylhwDTRG/F
vR718P9L92HG6gGSUpdJM15tKjLdpelikhLWgzE2q0nM+Z99eHl/pKZ0Gy4KRP7R1H+Tn1+NQGr7
fA+BjYo2Qz4/5GL8eatETQFThFqGOKqf5SKiVnUjTbLb9vzwzNS5OBz11p9nYM/r2UEaGzpJelcm
hKCZGhQOwyDdxSBAUb/v0akkfZgmzLGvuu4XD5RsP8PPgAfb7PMH8TcAVVtVXdw/dt4bWggpx52U
ChfAn8JIdDB/1STEfTFzYbSVyIJS/t8sQADb/+Ln/z4+ZTFk9XAjogaK9K9eoZJwMStTJbg21Bah
ZkBt9ZACesGWoF3oNgKKmT8NGt58SB+b7eIQsP8jbjwrOjnkS7wdRVToewUXIZRfTrujF14GIYGq
SNeO2NrreXyVLicisN4viahCtT7UV0O9PgyA7VyERoGm5n2CAbSgqv3tQVUXzAhXzbOABWH4Lq6A
aZyTC5PHIJfTPwvRRS9nfrKF6uzLy30Aaxy7xIUp6Zmd70tfD/SrOEjpeRMynYpGKYd0aWzPFDX4
evEtphj72uXfaKtD8o1XbmLZSIfSKUNXvjKff8KfKO2icEqDfqBqPNtrPfzDTNJ20HSdlXlan30c
ujKf0e726+pM5QSp4xhg6K08vjjJhftm9IqQitarlrJdPaLfvSzKBC1wYuAjgP44vVQvFtY24VzP
OpU7QkR+67hC40TlpaUMJaMOO6TvYkJygndq+JCMxS3VCDH4vbSs6t5kLFye/IafCeSZKrck8Cjc
pMYpXxmqNkp4mIt+sfHld3EWfOjd8aduU68LuNmT82wQwfi9muMs8KvkIYXt0A+3Cd8tQT/VplHj
emhknvuekl77LhzHkXsgLzYY9i9LCbM1Hsw/BxsWO17a/cdnPZ564fxH309BCenI7DMqdl9rjhfl
qnQfztKfTbASxpToqgA5rrQlHlpiGHmM9HFAEE6LgpFQdMO4nQfgXvhuL/dHqrOVT8djYyNrWvL1
jGV+bFJ5PwTHysCK5iox6MIiFPc5Csg52hLzNeEKnV83Py8W7sIN9N4xeoIv6RG1t6CErgC+SjRA
YylyUxpCi8TKHHUOWMMf9xixlYi/6/d3blTGk10XEFo29PtvRbNR5UFUhuw6gD9JrG3j8fB5pWEg
fP0n7GNsDfdi2q4cAloRPRqoYQi8nYmR51lnhRAecU0FsjI2Wlw4Gqrky2mJGNYEmnNDVsOdxScJ
6pvTJVEngXdY05fQo48ueF2qnhHBv2+ExcZZgO4ok9Tqog2YbqwoWl+B20BAG0o+C02dLsptrLxY
3OwEfgQHGfU1DFms/UTBXx+aSh0oaqj//moEQY9/ekZKT8gvHAH4agzXhVvJ6Y4aGyL5ENz6CkUW
S9wod3yJxrIwv0q4lgV7v93I1fF+spXjiIpCoUG5tnxiMVn0s33Yv/Ol60qkIzTczZ6Z5zoXbte5
wPnWXinOVldCMXy9yzUf2+comnLVPGJ4rx2Hwof194GcJwy7mbrG4R9wXy3G9OeezB4vSavAOHn4
9SwmbuP8RMcmcMh3rP0DYrAv/ZikVZ3+m8pnmGV1NmC7zBFFODOI0JBX/u49INbB9m+8d6zT8la/
PUhBBSHO3FClqKHCFlZb8826w/IhHXs5jzv0FY22Ut/WCCzvVq7ZVJiEP34AQNsNcRYYWiV7Keug
DX5UrD0L0l7u4TZ5jid/lSA4H27QrEWyQ0eIHPEen31hDr5w+nUC4iOnjciX5u0hCx0/KKlpj64f
8CdWCtdVro7VRiSbmDrx22bfW3FFeImpncy4mW2VnhGQa5d8g45zUlQY9vZ+mDIit/O7fWt64Y7n
mGygGfzIUTCAGyxAgYTb5+LwhHXk2BPEfhnwH7xSLEj8L/HUaHmjPL5dlrwwkyju5NZjgCTNpV/G
nJcpqGU50Y/so7ExLIqwW0hpjWLrBrO7kNPOD5RKQHWYiTf2vS3h7rNTuCuJv7K3/aU8qyj/pzoc
dpMxTNwHFzd3eoAPOzGFK30FWWc3r+XwiCvCLZYb8fdhbBTwVvqOxguZLzhil7EBjXmT1Amf3F3B
0k6EA1I6mpgCPSURyLfxVE94oky5qdOtx4xVqDivKE7MGXj/V9fwRCXcKboSvHcpNdeqBYqUtTMm
FuhPevWKsGuHMIk2BsimzU82VLZvI3ZLSZtYpzall6ylb3CK2TGHh/hrlLePeGXeN4w6Ev9ycYyI
IYItK5ZnB9CtPBwfZt4Q1tTdkfWd0alyB6PCGRu1zi4d+CzM+uuh45k+2Uknwph9XPW7hnO4d/CY
TcsqTopOEJhI87adA1oq4yjGed0iE8IFEnYLW1NwfLFPTVrh90xN/crfE8XV+OkfInmjHbtAUPZa
ZaU8XzCZRcXbJid0G81C69MZ+hE4RCBAoTIP+s4kPPN/hAx6jj3HC7Au9quzGS84ePVl6EXRozQ/
hQ8AUjw4k7oT7P63vfx1pxLQ4VzLckPishj52rj5KRet7yA8t+NAb8tBMreMcAT+hBXQEK/b1Ka2
pnumopYEbAoq5wXxwqqXuNas06Llo+wbatlUaaP/uEApsQkrvEshZtE0UCQhBJdCK8ZDkiUX/3ox
jYZCTG/sHY6mXHqHIzuUYsXXQCUXzhzVKw278dWVEQO+nOV+RL/PCJR51JLbksMuV38R3pjBh7A5
2eCdHieK+oXChJNkI+iUOkbkW2m1L7VtlDJfFclHW3XumeHlZpbU0wSSEMJE0fjAFohEcYLemL/j
P3pMtscrASEomAGEPt7/HVwY1hPwA05xBEQ9Rk/YMPhX2z26vuUiW8POW3cR9f+JC2tIP4J2/7eF
C5MvMpusKCQBrBM3xzayQY+0KRfqy6wyovB5phJpTColQtLkmcGa0y4kho/ruPXiGnZ7MeDBxPJR
OTEZDTkscQOg1JdjJ4x9uVTxo8ITQDqNCJqG9Hnq0AbypphcWAXeMXAWd2NGVsOaZjUXSC5UinTv
IjTiVT0k/g0WWsYJTy3UfMG4/7/bDeJ8wJ688c9ZUCK5PKAohg5JfKE8U83PO3/bKeViHiJOurlu
Rie7i7KVu9R8D8l1rXklmlwkp67YLtTsImjZukX3+9hGWyGYSi45Aydo7werxVJmvdo54bK7lh7l
eUxQ21aJtluJdoDtbCjKu5dV5MBgqEtP6onNgIiY1S3kZA/yUMe2TWbawdYk7uebs35KXhTKnidM
3hLIomNRyKRTcSEqUtBCk82dDYhN9K+f8JsQ2V2dmnPfGwlSGLXoVNwVTbF/xjgeMcEzvbZnN1ZR
TEwh07nugRqHm0vHDA+oMA+DRsbDDA3qHXmFHrlgum8jlORGHxV2ojLbrlXRumXJVrI/rx9pgdIl
++iqH5F9WqaYB0pm4oztKNyN8+BPWvF7PT19QKCnJ2p829nx7Ai/bK7nouPJdrMgIKkJOD8W9kgl
18011vfLRnagguADS9l3v9TtYtg6bv8Rv8IfgvrdYNo3FWr9xTjGfNpn2J+mLTZjZSKpBwxDrlTk
8J4DyRBIUDygcoyyKMWNWSx84434QfCbQjvvrJ0GTB8kigE0EWdrM40Rc1NYlMIGYU7I9lWz+9OH
PLrL/anYA/vw34KrnmPFPoZcNuY36usMvY0CjYQm1JHvp6ZooHva+wIvmPdYxSAOPhiM64Ud0lmC
DdYI74C3aVYHz7P1d/iC2SMajs//hxiS6RP8a1MSNKQ4znGhmrRTlC61VGMIV1jZR4nbEZ5DhY2u
WqiwOf/oRVcBjhEg1IrPTQ05LiSc7iaKZlnmX/MnWlS9PwxXRiwMvzn3laSO7PcraIM71ZMaOVQZ
yf0IEcN8oGB/J6qe52nfEFSrvz2Xtin2kCrtIPMcAZbuBPj2SUWsffErGVTkQmCKPUTTfBF4z1hL
Ab2ccY5wrfYbSTq3sYPyn8W57V8Ox+m5vNXErYrRgSvhnoq+fHgSpuGkzLz9hVQMeECGtrxJWgPs
RPQhWzVaCZ9VbEoi0E2clHnYWzl8NZ3lmPHkkUxrF6xFHgJaTB+eiwueyc/PjZBmNlNAuYPF7G7p
EIhJeLTD4sx9QF8dmXF8kF4d9c/YE+Lau0s9oKmcvdHtCGHuVP6I2mrPmxSfeFL86J9v9lYv73ob
0jrPwBxbkiKpHWYGnO1V24G1Nj8uJBo4jFjuzUs9JjsyhHrdNXerXgAXDHY9+gxYwhuZwNVQUeN5
NwtUOeQ7h9M6jK+7EQlIyNcO3SfoLI7Dt0JJrgYdF3iWJ4eekGmfK5Kpl9fswW0LgveUDubmrIMW
9ebTwowRPEq840fWtyQXbWeBzZ/gCb5UqBOxI78xIggbFJffbx0yegg9MFJ+vUfNdpsAhv01cv3E
M5ynaYoaIxcK9eyFn+OMio3bfyqUlc8JxZDEyFeanb98tb+cbozdEw/jqJTuB8Q9cNMcGima+EC2
cBYHcVZcZWB/By6PKMfhdC6X2HWVIIj1SywCC+B+lOqsN1RfSn3ossP8rR7qSsLLnXlB/VK6LFy9
ySrhHrffAe/RW+LNxthe9ellgatxvKOSFqChygaUGOpCtexFnSzsxrfNST3NF99j4qaYVUW72Ev8
kE/4SQL80yN87y/IoTSBFeCTUwPMmugreeZmNarJEx1rEY2XxMMmJ5fBtIc8I1YU+KVVbR2N+Fte
VKM1ocd3lYjO/avWlZiRCe4R0GpwKFBn/zRf8ZUbdTu2C1pmVnBXqtq1xKcLomO10vKYE06axnLJ
sZYE/JRlXuwTUr0KN+xPF3uUks+WAHTUnyyN10ylsZBobPh9VyBJejcuf4pB6AW3V1fneuJcQHEj
IH05jV9/USW0+b2gX0h+gVVTfZ07t4U/VCW2vwrMJSlYOy+oQWEuB0v1uRCkKikx7/1lRqMduRNi
2+HqGoJ0Ri817lMq2wCIlPeJLvw2O28T8bnSHEoW620Jro7bDVXuxvpeUEzlX7DHQIjRygykZAb3
NDbOB2cQLf8a+G6ILj0iPeMGHEyT/p55qBQJ1cljwb4daBUl9hHf0/c2JfDxlSdk+YhBGl3BYwGT
NjmtlZtxE5eyvNmhhG7Kb4rMk0XCN9Xz2Hez+/5l8a6lLiNnxo7Moe2kfVT75+1uGb/4XDQpT+tL
fFqhpxgmgnUPHKBKOI1eD33RBE7mXfdZMRDwLgYHmjc/CfpvKUAaBwbQ5Iw6SXAXcbzrYZXLSl3c
wKRTAUWNZV3nThxEJkBUItnsh49UyCeYBeAmkvq9p6ewn9K7QPk4pSxhFGhKZc1iauwyThJGIvZ6
/tKSEdeb8xVkPhJEwIAmHfmr+Z53txS7cdHJhoFxt8GC/mGbICfG5u7XJeqW+vUrfYog/khwwary
PwpR6UbdWsFTQC8655BBaiJpyIPEWMbJd0gmmqTFwq4fF1BvRx5MvpOULRqbgHeByU5bq47c3xrw
tiG8Ejcsq0ZrLS+Nd3nZyWcdvMiO31uP8CQ3JLvb90jgA90Z4W/iRlmmN1wQkDEio9nTWU9JJR7/
ncRO4zwCYkhOPB8VkliVRzjxCiYeUSae311kbQTX3J59qLUYSg0VjsCm+QstXUpcEvx0RGnVv0ca
+tiNvkUFAqxD5IrE0QvosobalslM7xn+1pm3RD8QHF9c0rDnQMayEBxFjaT2ABRUzMGbgWAUlDQv
fz9Ot2jRlpCvJv/TzxRuEFIZL3IleWh2tS1HleMDnSMZoE7lMlGXcnp3WER1Hz72bSrw8PCy35rw
H10puetBjHXgdnKgNAxocHtLsZ4ApH5BP2e730wRy58ba5lj4QBYv1Gxja5ElAKB4Fwd23gsNUYn
3az8sCQDDVBBM5m5P+GYym52ZYt8m23dO0o29JMqm7mtlTGUI0EmVr+/XIS1PFi2hhQzELIuw9m0
6BNz/PXA2Jw2DGUEp2sVNfmu8r3W7Uf41HUYsrnAOD8Pd4AcsFFQn7E5FfAL6w+mApSoRX9xiT86
Tkt9pEGGdgYCmfERXYTtx5jYYLYCxHEllrewS4pSYFyp9hogOKEfmC1v39G1pyBss+r/wN4SYJa0
alTkNYPMSD5XclM27ImDUiUhzPsn9a/KLZTWbPAkzKtx5knea0zra5xCxKyU/GqiuRS1VDAig9Gj
erhycKyX8hpL2Zx9ZTA5qrkXxAgCWIaLAzs0ALvoa+Ma1NSkbIf9wPxoMowz5TB5MSuyq/qKn0qI
8A571CFgoioGJv5U/nx/pP0QSqsBvzse6UbKehIQWcJB6cuW+FKkPEGQYtCk8PvekJzpSoIhj3KN
AYvW8YHp9xJ0ySiOOMgGYOgsFGYWrQ8GIToSxSy2VN5hdQjnYDApVMvD2sCOag40EIWiDQd1FW95
U7LogSE2pW2/kRWdIenGI0SEBe+AABCv5XzIxTfy+bdXA0AgCUmMsUhp7LcJPWgDR8QxJI1HyYr0
USWYcvBee2bibQVNFFLfE2qTmYaH31kN7INi5v2ZjRMMpYFBLue/NRUl95VpsdClVf6oTBIHhlnZ
sTgsR9/AvfQdEqqLrjHRWdCWDwLfIDo847PvmziYtqr63I1AsCTM9ZnipaKH+99ixPqxqTxDJ2BS
nyBvJCwmfUo9R3bpCCtFTipS+FeVAGV4l+QINox/UsbhUKxb6SRBDoXPYfzR0sUdWyMdS3/Oh4lw
dsgbzx0hCADk/1Og5X/BqCigK58TW2ahXoYgdslNWDhuqAzV1UqaoJZprCutMCEUbAgVMc6wbbYS
AG6rQLeGWcq3powU91ZgTEAitiKLh8NdLNLWEztIu9w7RhqkJdsZ0mxj8r9bvUDSjAd72WEkCiIS
KgTXvHB5WElDLZDEAJOjl082fUbFmJBVjlAqEGE818cn5j2jK5Dr+w2tkN2c1VriNUz0kPi27slB
UobS6NVNVXKsbORVIC8xO47yJc8L4O4fkm08w3ff0tRJlno+Y9XF8CiZvwltMXFW+rHT/814ZqZB
m+G4htRD6wK9Q8sHiFvX2luwAOJ7lMJoqfnDBuOctC0P/1xqKHDE7+U2oluNzmej8tGygCeZLgjs
8IHVw8Pn10b3I0LBHwhTkpBhlT8WQodY0Cg4S+CG+Ickm/zAnmJSvrplWSocNWNKPEcE8a5Y5ChR
tnUDSVHdpwMBMtUaNmcRBuPYy6JMqoksvC6O7aoWnz4CdeSnlrs+AgM2hfi4ztfgEly0gKyJ/flb
h21NER66pECqyuXX6660TGTN12QywsX8bfqTFoqaEsAUlM0Utc55VTD7mIcYnxW/P3pN/eO8Aj6b
KWel0V4IM6ae7FnfGwjShcZG7KMaTb+MyMf4GuhsUgaexCZzgwTx81ou4J6zhKA1YV4kFJdsZ9o6
NSFChYBVWikYyqakdeCpZ6mUd77QWQtRjvWCR0hmu90kTwliwRG1o+FAk3lG8IPWnBXaZongvupM
iLnbw8DEDDI6oY//rcliiBHiJee09bM868NHX2TeWy9c4bbXoxTtDNDV0mVeH29GnqNqYcrOjCXf
YTZfXd8gzYYFniN0iGxCaY7aWSKNhsFqVIwSEDEX5Znt0KXfBrTOVQw5TPsabsixz3KmHtUTNyfM
Hyv5CHbwLJI6gnnjt+DknVU6TjNyaD/pUvmYM8a7vmHgguy5j5tYDPgEDxVDaNaaJXr7PBbVOLcZ
1jdfYJHCRkQN1vdgy054K7XRC5+Afr+dp+g+wrGKAPHHNXQ7/SaUroHmsWO5ctOfAi3JyDY6c75J
kM/XxCptWHuWqqKr0uXCMAwn6Z0qTwRRoBgSFjY8N7qAJmz+mb8EInYHYx/M1enuEoYeHW+UZQTp
dX8ZL5S+W+3kpshnE2nZY6jk3dZYBTfpavR0rDNOjy6I8bkYhn+8bCdBTJvYRSjRmEYruhRmnIhu
NIateWw/Zra+sClFGQDVua5iXcsgun9ysd/OGwBpTnfTEF3Hkwe/cqpxxqJOWeruaqnmgLOGicjL
3cblkVtCVXGJ7N4etSV3By/ToUhLpVKmQyIOfv2ip1vHQefXHipNnl94u9KnfUpekapaJ/YLcLOa
mfNa5Ih6EiktqjOPjRRU+1WV28WVKH8aQr5KHkk5DAg0HU0U/YDDS+qbH8dZEDgWzVMmhj9uoztJ
i9/yXmLCqaDAJ+ctkpv5/EvRlIwnNqUwh0msPCPy7VaYiscuhP/kyy9fb5UIFj7I2hM03Bm2DAaY
O4+35RvmNcCZ3ofkYuduDY2TA3bbWh9eXUNjq4rBegMTxWu1JMthB+zp1hq6Mo3YkflV2woARies
GxG2q0FLtY9ogspu3z+p/5q0Sr4CieZvdm6FrGVoGb54HhsgoThnPL3fqxsOTIbf9Z80mPrT1/ZC
GA/I11/ANaii/LVlnIvhmGEjxfYtXa6VEHB7kx9vHWewmC/BUDqVcg9mQ0QEWwvPh0Ovis3TawXx
MWy9BcGyQKbaoqt0qcXw9R5CdyuIjsvHygm8TDt55R+CdVnObgkH3OJlFcNwdUafnVTilq5LQpqU
r+72ODV8KrhKM3N9JdfY4WKVtD8V/mFBm0Y7/+NyKBnmdbibLN1z+aQvFvdb5+WakUzYLTKnj9jA
EnYJMsZraRytSUpLapu4WV+kZEUvZRmufgINMhr9bjVrGFSHtlVTmLl8e4vF6XJdpHNTEdwfXiEB
UVFb0z/9ARUk0zVTOJYC4WLCMu8u0b14sfkl2sgeLrl4KiI+1HJGG30WsEZsDFEcj+qh1am7Kk96
Y5jUCGVyKeeoqWqVDYNRT4dCPD9gDFIC7ogOhuu7DaLgsku5dFWq03z4x/R0IM215S8Gp7nFN88p
u4kpGVfMpQmodcujS70AnPeT4eLzM800sduAEuwTsfK3VZZ7U5ws1hdvoxe7tStLsIVO91fQhpLR
FRG0tbVimiDelh7Kms+19MGYrxOhQ5ig16e296ZBC7kNCaL47pMrsAhU/nsO9mWQdObLAxO6DPr8
6cl3mdox7RpCLAz0AFolj8JnIkzY+p/4/LFgJrY80lrbIUJFa8/CFejH1hhTAEFRTkVglVQrod6P
DI+ZMifbFaiOURRMPbm0UQAAIp7Se/5x6cHJTl4vpkTXotMC4DFke3QA0SVsUCEqtg4l6iQEvYca
2BHXTvnCaFNgXPoCCzFL9Lh5rw6ahAdJmTBBl0wYCG49Vbjbk+ikhCyIdRUauO8L2hfKW7TTlOdI
kRQ2YoLqSDDmvd4kUhyL63jD90ce4HN4mNaLR6jfmJIERkTtP8FNwJeM/Un9K2rzz1k5tkuHr7ew
qpactarZW10XJ3MWV3hJiKI+em8lTkwK7UTBwLrgMhRA/BP0z+aVYwfcqAhzrqm2vxZKG/JUfcvZ
xapIhIsbOS10tGGp37QSDYT6GWFgv4FmGWgbGkAW/b63PLZkYa2oQtxL8r1yU4d7DWk6Pxej2WJ/
NlI3hKchYjaNeZ12Fif1uJ22bmMkRMNCNVqmxe38EPXRgQ/0ONR8jANNGnCLcOVZP29lR7/C9XVz
F+tBQZVamQF4ZQiRq6exdtm2jGfZgDMkJZ1y28vjiN3HC7OhGaN724Xp/PU/pllPm+DQXWqmnAjV
ExkYJIjDvo0Q5q9f0zlNVOKWOC72FiNkQEVRX7S8kR2n2vS60z8QhOAxa2WL60T2QgdBt1tXrL0c
aoqoJT7u/DGCOUI48oDsCWsEgv1Iw5vTGaDgYR4UJkDmqk6ahorvR6/ZUP7pvYHIoBlrCTS+R92t
sfapGDKKfeohT2O8y8Ai7i5vEJRCqiyV9mweuAHnJ276wgDQAgdZipF2zUP4Lw5udIJxieOEs6hN
ygQNIuxLL1LW2hNj/hOV9kPC/jd27I6CX9SwoBcYJjstQz86Of5w46wtzyi8AYEI+eo6XVtQPtJ0
jLlVJZ89WQ/fNvsieSCmriGoQsPFnh8OzIlCL9l6CLMan4P9Dd3kCRiqezpVRH7VplZBdgNbXxUW
rd37/N0Re7e7BaMGrKbALO5wydg+OT1jQXwqgflXevROFlMjjjBxpLDOJve0nrL1xwgKwjOxm86B
1a6j+HYV8p0Tr8YL1jOjyGTNw3JR5KolY0eFhKz7EncZQy1HPPy7KYM8404JwHUY40C5J55lQ6dy
9CCaN3fAazxxr7ISM+7QJmkaqKly7ViniCU2E9+DEUXmjDoMyx8HFm4X8f5Q/QTtXObjmjLZgcq7
ayZN8Q/PjXrL2WvfX/cJVsZSMja+845uljvMtuzIzf8usvGieSiQlRjdwUstONxVM7wj73qjDPz7
t0fVDrgIBfFu9VXlyPU7Umscd/QSh9AotPJZg4J57qn37enGXhE6h/1OxKxPSDc6bSo6zphepACH
1Ng1UH3COySK60mkatcE9t8zKIJbYlC0MBBG0PNkAHW3qmF3jwUyHD1NkZ3T12nGV8ZgGGA90p8v
4xaud8coT7BDGJ4vwEdpEYO/iFae4/+ZWODmaLQqxPHZoAY1VJLUQVr38y3O0cbPbWjIeCk3FgRm
BTvUyq9qHD9ThNJZXHz8Nz5SWRzMrQxQjpZYBhxyUSHA4f9f0mj1I7eoEyrDZ/sravXht+OiW/dz
qClg+rLn08xRWTU+0xR93+qi/Rd1tKt1BqQRQRgzfH6xuEA9x1OZngl09Af2KEz/BeDMZO8BIcKL
EGuF6Fjtgbw1vayhOemofr+6qfTby7Bx86uzreylv9OqWMKIX785R6SlqT0N86J8eX2qc1E6SjWx
NexIqtfQtBQ+TCxrtW98lreTNPRTD79ThTwrXsYT++GaTUZn1ZEBjwNWQv58CD0jBi/1wHCKOzel
0YFi98zOYFirZ57DQ3zXiQ2oI3hqqaH+kaOvL/h/SaSarcGCnzgW072JW21Tl1ybNzs6dmyR4BDR
BjH0OJVvjK4FuoXXwZXtKvhygpHQ+QO4ujNU+CYWVG3y6SpDj0ULiZLzGrJU82osGz1NXe9Cz/lk
P1vI4PpOrhXs7Jh/aHQcinI9bIU4Gxi+eJVp5JDIUpltsdBWsqbG0rtYr6d+gz/ludR9jFWCSjE6
gMFOD7jixsTYh+IUnTVh1Xs6GI6FysTP4bKiCsP3XKjHqYKEuy6s67wwz+ZStSxYO2hGnWFSIk8T
mRrJTz+TnRN0GJXhlBSpFBbQr9WQADhqsBhEaUFgmu5HK7LqgJdQf6L3LHlHMcUvU2CTFAdWdxKG
LEr0ZsLJMsOmYYPhAxrbavvSzeNz/3ffO+IGn/MAcV3NMDsBIEcSU+cSL9neZB29vYH94uKngfQh
kSljIc0o+jJCfPQGb+0zwLFo0r76qxod52eZDWeOyRwhnI9wgJawsgZHbgPO5mN/NWCNYIbJc2t4
tPVo6qk/RbUnHjnZPt7tT2WjxjzqNl0kyUVuCQ9TWq9W+0IbkXEl0pEa4EHqUZ7cI6HED2J0UN1y
LvFBKNMd5CxvXuGRn3fg68RvoMN8StOFzGDRM88PtZ0+/IhQYm08ExNSS5UG+TqcispT+4YnCGfP
w5epEIZYHjCxEXGrzHxiuBEhQSaYuhWI4wmFUyIN0nSB/hSyLU6IN5Tp4SJhRnws95SQbqY4y3jH
3Zyc6ALdeP4bVlhm2EvMNqv3KnJ/fCpLi/szKx5f5YZNKKSuu/r9yH/QyOfiShBlXTC2tk5SEq9N
Kn6/CvY64RcaDkR78e7PYB7aGHgwMpDxzFTryhKCo+o3xsJQJyWYd/wj/9mIfr4aqp5k+DZYcUZ/
jjCjnUT0Od8ABu1Xh8WnU9Y8CD1lNu/QiL4s02LjirLz+giO3PUTnrWbT51FjGIwEXvVLzXD8peW
Z6WzodcjjAkwImczRGV8nOZA8CGvOQTYC0fOhRb7n0zrE2/UpEZIamsITCD0Uk8llqSMrc4Ui+Nq
zkJUAbQrzYsP7fL3Iqw5A6GWaO/MGFAlKqSQ7E4qE9FUTYFL/iM2w5bO7GR+uxEAPhp03cEx+uZt
tlxUZuoX6foRRdUu41VIUMuk3gx5ol6JN9YatjdwJVqrcROt8SV8dxN1ysogiGZ+vPFpxjetV49V
ZegU0rAaviH9jNy6sWmKNC+YEySoUU/+tTYXt+HmVzfynu+o/1Ix9zsDcT8VR5f2tckUqlebWFAL
zyQo7pveS7+zGMThpb+qouWjTiSK5pkL9mDgpHuCwOUiiiFKc+0BRM/XkZOtHqDtt1QCB/jbQKxT
R2ZLZELxCivP/XiK0Vq2j3Om4I8H1h6+GnDvHL9JzbF/6aE7+xVc+d2L5w3hswsWh1qSv9Dr04Sf
v74iRtpTXzJn3E7ulUiLUNWOQN/JUBoDEuMPCxXVadF0gvLH299JfnBOSQ4eXtSGZJYPmHbsjp0O
BI671KWnikAUQ+VhSIcf3IuR7JJWXP0RRIAsD8bDlpCJgzl0weHMc93MTK+TdNle8MuS7571M8L9
lO/YWCeb7Ss7xKjt09LwaLlE8PpVWAn+bq+mrKBRo5LhTttEGK1vbj59hmBK6rzf7O2pReBLTSxn
xSKuRKUwZtUFW6z6sBdMYUU+f2vaCkal4PSPyJSwMPLfhoyKf8kSHfQZN1NHqA3F5wsaoWYVm9af
Mx49e+C3QqkA4sl0yWZmvX8rtwlpJG72L1m/bEmph+87lOZiFynT+QVLDxP8kIGDibBbXGCcFeFO
86tV/rro5W6cF9tuf4yMTluRm5QNzIK3/Bg9IsepCuzcTOkMW0JzzDBIBkQRuWdPkP8Cq9b0TWhs
nwQ1wE6K4N6TNfdbc0LYlQHR0zEVBQ7R4LAcaLi3k6LHDHklcOypX8rZYizBBd7c+IgPQf1zvLoN
x5vqj5q+2kIerlDw9SL0uclacEEJYgSrOVUNOjEuDW97bcyGp59w3o5vuJgOKOe4WtkvaB+HNjjz
DNghBzL6VsLOIL46rSoE3V1pokq+UvcPBLuSyxT/UFKDsbYWa8dUTJDm7jo8VwU9qulTtRCegmzM
+nazTjPRxSKTgNOKcsiTXYa3d6jYP48TNIzK1QP89NixHVerh3Da1drleJDJtXl1J45DQiuD9mqT
/2v8jXOaE5MEBJCvTAtmI/L3BYVVqzibLF97i0IPC5CJagGnpWKO9Zq9GCZYIQ8d9Iy14yVM6v1j
XFpPHxEs9XTmJLHiyWqdD2nTQSvsR3TIns+76kF9FH05J0h00bCB1nS4LN8pGtdmfohAp0qrzjYU
10rJFvfBJA9sxgjf0p4o0mRx06OSVNP6xi58MLYsFjiXpaKMpM5JC/nY4LiMlrdm1Ltek3Eg6u9p
n2tjsakD2VCGqqNgeAjh0fEKgXRH6OjJEcqHZsmdYqVoermS8MURcmJmXYmpIdtChrLPKaKdm/Yn
W9Jv0z0RJ9zgdKPDko+RoqYwQFVZyYGBc8puZEiy/gBXhCT+ySv5UVl7LeBcQPMTMrpnbmhVo/Z6
h2g+tMzvBv/IQlaRXlI0Z4MP8C3QVTymhZzKsxS68loR3WOq83QCXqOMy6kHXC+uFN1QfOIrio//
hzF3wLYZdeiClnnmo7mQeXuGeW2iK9AL40/bjFWO5M8x4nJ0E5cGySMkcEbbysdACYp7if+KjSKJ
NPAy6sZ0/ab0LT/YtiE/bl/GWlxWH+vaxxI53IoAP62MumnDdeivPcgcVtbBLbT6bXBR6J9ci3go
OzPApEJwd72ujPw3apAS87l4s7nfF/0kz5qyB4eWlC7kcybc7FerEbY/rvi/72SNSIQHweiv8Va3
TZh5alBX1vhcpVi8hNuv+Gq3TPL5un7DTgkj50wvvYJVP6j0ymvnoYXxnWIJKMHyDE04ViSTWcBy
KDcq4/s8pa3PzWDzaLYim2sxj3+GTgTviKEjvhqvrYuQstuFQpCsvMpqh6Q67o2lFyAGQsm6oSfl
/sEepTA5WNqZyrW2xc9owHRmw/dRAS6TANqWPAe6rm0C+/4tAed4r/GeKmtxy2FNaB2w2TphpM0p
qkrlu+aCvDwy3WuSBrgyBAS4+KbcRJUS9bbc+0JSTxCeCQh56EtfAEntat9QiR1ZR+/I9Gb6U+oQ
NS2Ay0izKnRjp3YXKd9t0n87E3X2kPFTQQWXXTSj+nbNkUBqW5v6QLog/couCo5ZBCj2E5/Pmm+F
TyPsxjSr3EB634u6qPYmzs9ULD1BDpHqwMhkNmOHRD8cRX9b7/39yTxiTwv2KwSS9FDWP/Q7+sEl
x0kqG8eihTcJhDYAClEN6IUPusoFdh/zOv6GmnRXsGtFDuWAKB0AVMgOdvDbqMD+9ty57wQ4j1yg
6zqF2tMp+M07ZA8KBeSPx7TuMa+8tJRY03M+8epOjKnYynlsi3/fyg+P4a5jLoZIPMpLA+azcegQ
zzFbioRrRHChlO/Qrd6TvAqdhgbl3Bxvnt9tlR4sK4bOoVAlYCtoKISa1m4b9b0tCypNx3XW/Qby
3AYlz5bshyuIpALjM8YdtHgZRK5ZnM3Ez/JNiq5/K1jNnkeGOV1mH2RWFvPcz9EqlyYDRj5Q+kiC
/RzxIyN+UA9AlCZu3DxPeYwlPtunlkG3mNQdqablThlgT60/EjU33Hzjm9+6kaUoaemMpPOl3rKI
ONd6TbVwNnsGsrXM3BvXsASEouHOEToGrn/6ze6NtKiV1qREvmnVJPz0h5edzhsJ0mKJfvOyDdjI
BkgHF0pkpfvIrbmnBfcDPJTQcOkNmAOXeqEp0FHlgaDhMIQnn0STOy0KxVxkNuk+bFeWHMufNt6B
pdEEQptNX91B7BMPTzoRwUyG2hDL/u9nZDO5FfMOsO+vWBLhDaVvO6jy0/4XJeK8cxl7FbAnpBDw
HWYjmb+usOFQbRpk1l41D1yqOVs2Cz2EHDIE89zxDktjHQo7uNcBbKXtjSwgxjTwLw5755KQRG6a
3TcUAkgYiQfzU21RMnszpu2j7hjWhVLIh5JPdh76E1WzqJSFCRnxfdisppwFCHJYhFuweJxnq9AQ
gCqA34WPeq6J4tOuGgB5/4H0toj8+0EfsgWpUIZ/XFVK+gysQ8M22YlWmtSf6xaX76aGKMR/mIkq
0o6BBMruB7x5ZcKjXiNcO1N7UsoSY+b53lasJF5ZskG6dEvzy5KMwhg6jtZmIWCQ/mm6y9cGrms7
E9POeGbP1eAUGg+1+r0fblWJycbcwxi3FpBUUE6qtKKNMx5lNxZSZ3ToHYcLrd3poFQsib0vwNR8
ixcTRV+TucQ5C1ElH1hEb5SRAQkHBjaG4q35itTND+aLOlP1epw07+V83jCgV66yqUMicQdG805z
hjQlcV+tprBHbgX5Pe2/U+Na7XgVEobAbVNob6ogdjAsIP9RhSECgd2CTZ1cXic1VNZ7plnhEGYu
3vFtLUZ9HADPY/Mt0I3DpQRYuo/xUR2RS2YSl+EyeyDrN2mwF4QXseivrjzNWP4za0RUrYNwsq2V
rW0qkwLboqtzwQJnNLvDB+BwgmsroW1VLiUf2yb5xxRSjogF4tU5uHr4qNnR8hZ+JHbzG3uUuenD
fyT7+QmAgbkdzPrtZtYhUwih9l8mHP10r5zVE/X6kBtPfrX3hOHd7LjZXXQcWnEqmG+5PsrGU/dq
Gf2exjJj34d7nbxrKtw5cuFjGmzu+l1HJ7/PyxMz+ulquSVLB6W14BHHesdyH+uBq8qdtO0pAla9
kWxIixkuzVuPpJzqv3NEDjxT0h6XMG0mM8zpwKddppPSNtTOByXFR5FuPB9tHIbB9MKnbWZCqwRi
kbS3K5LyvuxjWMBeH36O5JJeofhUoLOCnARc5jmkQN1VUqceMCyujV7Hju5ZLedOowSloAFNk4EX
LUHanql1rQuKV2j1E70ZGPxyUw8WUsEq1G3geua5rLijN+ZUeJ/msGkadAkOUk2WIuwnyIvs1Tie
aZWFKuyVxxr1+AbPln25uzRONq4oTY9sSL+Qd24ynE11aR5RPBgtxZUKsjkva2HjRqX5QexXSUjW
Xwll3W+kMgMQDKqJOX7uAufz0DfsdDamTaU7d+MU4+phVBU+G20sN20zFS+jB6OgDMXmEwrzJUGh
NvwFC2AF9+fybnwHLnhljptB9SOOi7GlpAC/g56XFI5Fy8KblA94XveDnndwUmJY7coWS5WP4XH4
76WLjn/Kdx4FVJ19O4xknCadcgL9zRj2pGtqJkcS5/0nWCZUpASXJw9yUWBeDY1D3WM+LksuE0u1
qq8UPQkJqVoXOwiOgkuKBGAC0r5Me2dh7fUWrs9lkZzDDcvtfVso2h+c0uD0x3sUy+LkFTNTHgKI
l1wKzrK8PXwKFkopUvjW2DQpnX7qx0QVURoCeewtd3b+bDNSjP/fTfWGEZuwWwIxsv+m+oe9HL1D
wGwP+99m1i2VWkbbxsGRALdAU0BEUyDdbJP31HYrwhE5Qo6m7TUt//sXyO16n8+pd/BJRdKymM38
kH4o30g57nmZxfetCCYe+JEoIyUnACD42BUjH5CwME8FH5NTHhBs6wjTXo4iGlMxASwLsSUEjB28
1D0Ly5VJG1aylq4bquzJnB4mxEGsxACFCZqg1ZauzrtDr7qpO7Wltfmp663nCpKIfY6D55b6s8av
OVyjI6nn3nukbalVOP+YeTLeKxG20/nvtTJJopCFVIsu4HqoJKjiFFP4gEX0aYDNgZx7DarYRG2V
II0nMTY3CjMpjz7By4CvDVsdNyUuKKzbUmwiuzh3lG7j+LYJv9tU/fO1VHfP+AqSK7iMCVShIa3n
QyNPPMgEkawkcsuaenabumXiZ4tdR8nmVFz6WLlpHGAM3Vd0MYDSOPRkXnXFt7l0E1pHABD+YnVN
yPblZqArDggDUvcelGdcfDFzIHZi4FwoEG3gBHwJdj1cFY/dQQtu9ov7+nzPtmKvW+QBc3wCqVAT
p/Ew/uzIuC7WFCfA5EbWHnOlEzEH0UgkXH9ULOgV9GnH1Dop19UqeuzJ8oQg9qVD5xTZBOtYLrw6
0dtuExGefW9XrmTK4JaUAWUn98J1SnNUgiwYojR41eZjc7zunNbM6MO9pI+RWrfOLSqJ1eRSG6BR
l28gf/8lIdKyx7ZJtJlboQ7iTxkCs6IhUrdk6HC/f4jHsVPqQg5AvVrxxcvaC7bhEbb5hLnuII/Y
55wyQaM+PjrAC8spOGkyMP5CJ0vyv5CoqIGEypwGwROKANORZTnuX9Iga7h2tRtw7kiXoCHiGsxJ
9myw9wchrzdc41gjv56W9lqgY8u7Aasd5/4un3Ga0wrZum31MZIMDPTBTyhT1GpDIX2YeO5siMfA
vgOH8LgWzgYNmQDi1ETdVfHBWAAlC8HCCCb3KGgZSN2xwXjtH+K+Pmem4geHKIQwrEmwBmRYeY99
ncBQi0iUIDUpA2KdpLGh/u0YmGywITJIO28qVEOA2sQFj0EaMcaMU1KW/8/3UlRs2RhUNyHR30x7
pSofq59Caqbo0Wg/+jFoz0xo8Q3caYPZ6fN83aHgKvDLiNmT0PITVcNxY3y6/qx0JOkNGqtoPu4I
N58xHctTtU8DkQ0G5wei3cr+ysQMjbmzvIoIrXbxIdxaJUhWns8VhkKtf8oh4LQkCjpCQ38sZ5yP
joXqDnPHDFSwPVV1KpMvbi4wT6DyGjN62w8a+ls06Txlcf9z1YUDQjP58Fn4ofDePs/18lOnFyaq
xGg+wpq8oS+I+Goapbm/WrdEfTjYLv3tLiy+SqNvQUiyD7vRcxwBALbWRQDunTv6kMuxUd2YgyP2
LznBAzIu2rnzO8TcTMfv5jae13XHmJVT+3uZh3bjPUzXh9I2p8TDRZ/C4iamYxF9a2sIyXnmCpo4
aejTSIvBBdaXGVf6dExVZNi0MlK7zavtMVRTyAJdXqtshfdGX2K9zZYRUWGPaSi4CQBg/uUVFRCv
GMf+RhYvyU3MOeDKuWjWtRXXTq91gRJpnyHG8jxpz6AnWwFelUVw8l4s1GPVRQ8e0u7NX8V19kJA
cNnuneTdbkqdwN0xYtpIQ5D4+bP8RbbVuaIoHy8DEovhQrswBVnPS18kg4XV5TYhlXhFDRaa4ZkC
XnXcWfb1MaIu7vel1PYNDjAZ1x48Nnk7Uj/RacutveJz2SE13HgxMUUG0Fh5K/YMLCbROeMzeLox
oqvKkxudoxrn+WtreTXeg0LiNpjzn+k9XTIwJunYdjJd45Uojg4qQoPahbGnqyLvLVyrrBQuvq/E
YOu4UVc/o9Hh1smPLQYECa3Mil7hmpsCQr58x/cKULbDHc3qr26e8rDq4BUxlczR8bIFid/wCaDU
plgOeU9kdc9Cwf1gZcU6k9A/EhwA0QZARG4XS8A+umyITebhv+/fPUyzE7aliL6y66kVZ/9HO/zZ
ZZeE0uRlo/axGoKxvPaqVaLrWO375uyi1l06EHr4+xLE5Lcj7+6dqXEdpdUhNAwaski7pbk7XTGI
SAq/Gp2TqCai8B/hh8UC7etgxrkQpysmmwD4PvQe7bnKp4BLK+yH8EUhRcwzD+FX3YzE3AcCVT/p
l5+wwuNhjde8RqpTQauEY9YpyzSFJUJo3wn+HAW+BQsjAKka5RRHyQEll7rlns7EOwsQISyrTWSW
qAEoymWrGqyPgT2YY+cBmRpJcNzxAZYIMarnQiPig9F5v9Jf851BSRR4hBwHrPQAxYfrsauZI23Z
kq8Unf9rXVW7ib3baNVH4qN1KUexiMgPsqNX5x65Wo0uXD0d0YPC4qhw7x/A7TGvqToCN1wFwucA
fdYIuxhaKAjy8yLA7QvyWNR6ah6wItIqUUpKai8ohdp+6V85vSCsLeJagZp/vANJ+IbrovEaM0GG
ylNWk/FrTMO9BbMcT5Y7VtCWX/zHOwfun88tk9ATeaJNnJv86ryOUbmxQPzYwXehLmrJd1v8y5Cs
w5bX2jKXuQgv7Iv2lB0AseUuhhm9c4hR9fvjVP96umffWM6x5DbDGiPr9298hc6pzGODHOfCFYNo
O7Ao/+0Pz294LW5UXqJMlPgYlUUle/qS2/qztMTRDjjsnTcCbCBRrGpwNlcWkbruPwbDk/ZuV9o9
vw7PG6MuG6LnFumCZwkjYiSz2HcImR8hP9ex+roZNe6EaKvNn86Uxd7cXauFL/5JWTwSQ+fG7G5+
P3EMd4Wii+g5Jyc1+2PQdi9Vla3zWMG06thfr6Xk/wbVFt6aHXJhLnL139z8OQzhw+oIlSjtb2Q6
viKFTFVpQwVURT4f4hQXqxgBV0oiywGw20pX8mUaF4L9jXuSKO7ZFjyjUP/1oc87n5wUD4JOVMrh
rEKvhT60Nz601ow0XyHfPEJWxfie6trlurRajxZavWZMkfNiNWQLYLlqTY7M7hSaWXSunUv7pzj8
If1IkuIRHuF5S1H9SKmAAxiXXLM7G0YR1GEd+XomVHPg5uMA7CPqenQy6qz7MbcdhMnptjjLBoZe
nZzWswDmuyio4oqIznutW2Wxe4NIRqksc1fptoHPwl11s9YxMjMA0sP1PXRuhK84LigRChlnoJjf
fZOfidwhppGgqk//YR/wJ2V4qzjauSVe8CAtgU6fBF9X3w+HgQAvw7kqyi+uqfKNm8PQGoZkwLvC
s5vS3pY6RXwfkAlS6nId5pgha3kOmXt+I6MEPRbSku59vQCPokJ5i3cjKeMFgE6iVmXWdjoIIAro
l6KZsoalxzGE8p9S6Fn667RS7uWcb/fCmPxS3Zy6fluiAI+j7+N2PFGPTGpMlw6Sq27y1gi9lrNX
f/xsmSrmqlOuMhc9T+MnntQR4FT1kyXEchvYvrszfIaae+rTp1sLFM+D9Gz5r5aasDbsg2otLCuy
ozYdHeWQG3bbKVn5LDd5RT6tEvWkQmikaY22ENCiVeLATz4D50Eq/uIgATMYMlLSoEwCIRoUitNX
ctt1T4Wvqtwa1fpdb9g4gRcdDWtVWWlr2wt1ql1RizCewW4yewphnKQFXao18gejBgCKtLnMUc83
m109mTM/Ii8g0t9hiu+b+FkPE9lS76cD7csO7oMirtkuKrpuYFhypXUDzyHTRRFJ3p8wP5NWUmU6
f3Q7WAjhf0M9fts+J7klqqViOnxymTCW2S8ZdTlHQGiNuaVFmXBx9oGSXlOlO0jeepUiFROJG4dO
PhFjKd1tqzjRkhK0PvWtailYndNr8MRqKQSLOKHZpXrVGNfc6AfAYwtunZVnMkOZ8L1alA2+53LJ
UK7GAYuCDndF20oanGD3SVxsI0ZImLr5cqtGdYLMx8IXKM07AZn0FWkzKJM6t9Tl3D2mTfGMh/Rf
fzDTGEjSHc+7Ss3N0/v5DcZsJtTkqV3BtKE+7r7VPMx2bVIcgO5VVD+Coy5X0ZXJX+VeUTXHOAuI
Ecl9VQGpwN6wt1T57bbpMQALx5LK7n519gh4g7ckCB5DpHqtS9tTxsAuhMNl17DEuF4eTUYkGN79
joBm5pR6+k06DLhyE4ZUlCzcY5sOOkmaL1mPZ7gfBy2JMfVZi+qikbF0+MTHkQNv9+HcO5zCIqPS
a6DN09hnm7Qw6kYLDUpHv96YO1FE+ptPCJLCnFjCOYe9s3MITRZiSwE/A0gxd0EEKHobbjYlvg6w
i+YTa6XxJ/eVme0GAxM8GdEZKw4GpXPVE5i9pjftuT2oh5Eutl7poVYt+SkvVDoEXYlE99zANI9y
Qq788yjuBo1Im8LimY+TisRbvQJaCuq/6mHYZApNUO5dNrlJH3n4paFIoocBDvsGF6UvUD6CvRLM
/NzFvq/tTjZTIXRm1b7PTPIqzikVdjuVxRSIuRErjNBFf3MIViwr4LWy2tnSM9gEILEcwiq9Howe
uWtb5NOGuv/ZeBt81KoAh+HXCFAvXzj53McF/WpgNiYf9w6UEmzBkfFotYBEzFSe4UelbosSCHzx
wuXpaCRYuBOlx0AI3TiLd2UnJywdrlyantnU/agp6RrVZm8PVyES2kHcxe5NKBjXVM0xHN5r6UmJ
WjAjBtM8r4E9aUgb5KhNw+bglHcIPaTlj10rYiI4ZyTQY3ZfS1zQylDw3CWWXRJq0y24bit+Kx0q
ejL4o0FgY6RKYB7RLOB46QXbu5npT439fqyV5rXDrfy1oUtpHLn7Za17BJ9YmcUY2itLrBt0LzPS
HXCdakayLf1RJ1tp5a8gB+7vJXgv6FXQeOhqBV2av8t5I5gACswepMA1/f24X8PER1PyPsAvXgHu
752m/LcbGcBy0D8kZq4kbUnXuNCvRiABxVlhu+iaAqD1Q+f+9kBp/NGEz+BU3m6dSTFhttThSYxk
VJ+lRmd00RUofJyg3N//VsUoMQPEGDuajca6lBgeeAYvVajKd8Ap2wtZujrELuD7gPHAPQg72TB8
54Ztu5dFoY/RN3s+j2DxVhc/gnRFlhtRsjWdgkQwU0yuTsXJFwoUr9GEUJe1HyiGqBoCbH33FG07
Vx6F3I39AsfUHQLlfebN//AsS1uUOmxq2o0eZdYPem7Dton/Yh2hs6LHh4ajckepvy0gxaQNya6/
pUoVHRvUHXPApHl3Z99O7grQni/UtjH5fjTSqD9Oxr+jQVUh6CdB5ym1X8d3U14Tq+tgRvUIOS+m
xz6E6J6RkywUNPQWUt/2l0fPPEaGhlEaJswSOwHscfxQ2yIIEzS98N+kX/0ndQEDPfhDdGKJmFhe
m+tsrdB33Osuqd0L+m/9rQvUsG+rfFOroy85DhCEotFzB9GaJJ0uVO3kXms/QIBbMakHqtnUx0nd
CkCzPV7bZMguAfcKF1yiveWsZkDrm6SkQCZB1KfuA6g1HSH9cMKUkHmnUYfpfrTXr2r60JuvJIV0
vAFQPDbWPmhRXcEg09JvOQhwIKymXu3K3ZW8KBoUnI5bXJZUW8cL5JGFkq93tfWCYi/rESo8ft4C
o7DbCFObL1dhmgNYvFbn2p//EiZOJwW/FYL5FM7PfIr+sPuYrNLHJIiXjJrFt80NVH/Vwf5CIaoR
BNPC/Bv6hc7h+OF9OXek2qHycWJEQywl59s5TEZ6JE/pmIfdfDBCUVGxNIda5s12pUCvDiWon/3g
8xfQrBd3x9NmwcIaqur8B8M5ytrOkOV0iyDowkpTLXS3H68ScljBmKGA5aPDwOa3d7WK73N6fckz
TJbdOSO7wWXp867p6n7eUTJHlnDLH36DAZ5XLBdiQYMI/aaCIr2ezlxXuk4vg9ecIqiZ9JA/rss6
54iPdDN/2Bj/yV1c9kMiqJcoaeWNI0AvUTAxy0yZdGE7SMpKLoZa9kI+wjLxSTf05r87BM3G2Vrg
38rkMAfgwxhrSyvfDkfvGE6Lcl/IQfLfwd9uHPw7BpMOH6fWxdFNbV6mNWpgC+Cfxi8e/yd5YJcg
/lF1qA4GyuWQW8IURf9xMxvr0xP+um3CeFb1xtIVmY9iehkkKLBWuNJoAYDWLJuGm3g+DnF6U2PJ
LD8Ed9FdwANwLIQtSAj/FWxYum6XlcTdtVbPL4OyjnhQuilIkrl5cbphKC+MYLeMUVwr5opa4yt+
VbNGywPDP9eGFETogZ3h+wWJRdGR3cVFllNfIvY3OTCPYS60tBQ4RPD2ILDLFU6o71vBPUxF70mw
2OPLO9C+rWQyLIyitqEhO3RVIXr12KkUzE1/ZCxfrtEBvgrXejWByImoBhnxa4KM+QgxLnlEPJ4a
NwQGeTXzqgfe+WU8xUwE4Y0gywZRhIEzpVpHnCZfspYWVMy/DvKaigF+yZXfMiCZJ+zZON6WkwL+
tuYaWE5bQesoo1Za8BubFw2YHSivdf2YKUYNvHtvm8udLkCiMNoK1wy0QzoHIx1Sh9QgaPIzutHd
+3CRr26h6UjYDDaGMBTXHWXDCFHqFoipKmy2paBY3afbU1Ul6/pOYPWEoCSvVdw+l1ku712H3DVR
zy1rsQpGQNAELqJequnebX4trPgGdbjkY2m6YfdRRUQ/jN53mpf5v53BWMAFdyqeRk/RLOtjbIob
IkEIh5fI8IXumd1IxUm7N9t7Jc+I0Tl33mBg0Ez8g5MKgZ4SoFgCWejJQO/xIWqlDL5SbpwIuazg
8YLI4VAhdLKgpKdSycHVDN+LeOFZ3lqDQ4p2EYD8EwwE+LPbgaOb0DiJZavO3criI2gCWno7AI+7
m014JM5I1Okl49iQWRpusa368rixpisCT38HqR4GqZs3XV6gTu/oNKJ5Y3hOCw+ofI1REO0QoPKQ
dVkgMwOqlJHXP/c2u2qrOuYmSK1AvALDPOZhvhxJ+e2+F7YCwYJfZsfoQZHwDAFaDRF6AFJIUZY3
aaDnWUfsGHuN7mKnigzI0C+8KQVtxZqmCOgd9FkSQpAjZ9jkkGJ6mGSBMcRiQ59+G1pwmuTSViUH
Eza0tCRiDBi69GmqO4cmJGEXMnnj9fLhT4k83t4ceAoIPQjfR7QBZLkBIQm061Snws1T40xiakHk
fqTB28TbeTfl5N4AztB7Pix734to2xzkiSYrxTvMEN1Xkct3UD0W485dp2VHTdPcNlJVfDwveR2U
XgfvTw4P+EnoUzORKjuG1Qf9g97sbm7YsAukxfXPMhEnrQFamfswg9VILax4veQJMKps/EgmVC2C
K43hLjWfWpg/yML2WuO2ZAesFAbjEzxbJDz3YRnuDKQLEHai1z97D2/s/xEXlRw0BA10bEOm+sx4
C9qVZj+BGPAgVdKVBK0AROPDFx8KwaRMIx9fYIY4VtRc1a5DjcAoX+m9/UkIKvgTcfWSskpR5voX
8bM0jsqSViRqF6S0LBc6/rEmxbsztmZ5MCCbRgHW8WxS2TP7itZ01QTy7fBd2cizhuS6QmOtaMbA
cCYe8NREGPHjpX7oUHnISFCuizusTnF5Cr0pYgq3t1yzxZ0v20rDltCrsibJBNvGhRhrVJ4RBsjK
d8FSWTkQ/dUmTbD3S0kYsccX1EtAE17ITYrTM5F57vyYQj9F5/RRT6bZnScPAmohZju+PxvANXAS
53AGSbCrwdYOhjBYk82UNEQyHBMZRpxmaG65pFyjpSQ2czTMJJv7fHVMG7lW70ZCCdTGuFQr3OG4
sNlZz75HSdap5jAmE63jEdmsQsnjFhe5cZm5jYy/rXHn1pXZq6UHS0FY73huyl06e54L6pe7pQYJ
+HsJ7DzPvEjsPKNJTZpdbT+BM4LUDOYobUf6MVa0csT2Fnwc1ywCrAd/a1mVpzkYQtTvFweekLS7
5kHYne3APPXyOrKSDDR07mRLLCl8UzTTqJDzicBrGPuR5ZOR65PaOdmGwH8rC7wetmGKy9kGb8fQ
uz/35ZSzEFYd1rm7WmIS8Qzgn4BrOCaz4dc7MzE7ZcDDT7/EzPhvtVABSdkWJCchzT81R5drIb6Y
O8mGEVTyCFoGO+FBAVexia+E/SYO7Jf+KSnCxAu6LzRto8oFYag+L+Viq6Y1t1w3S/HLwKq7yZMT
oFhaPyCWBhNAW/6HJzBQCwbCcC/7nnyWXO/K1SROPfgANVnf+zS1l0EW5B6iHOTIdb4i6SusL+j1
UgLcgW3UNWuzSrX4cIZ3GHX+c93ykPyBSAjySOilIznBCw7MCDQaMERgnO0QIgjBqXBthy2ZOVCY
2P7BgJdd9HTl94+IKeMI87MtvlXppn6yaR4UuwG/Ojhqh4ybY6JHe7O0Fo8EKa6BWlAcHGr+qzsf
wgWQ6I7WoebwWRXJ7wNgQ52vIPNQ+h369mGx/NJ9/1a319wPb8Mkd5IXU76qK0q32bTMH/CUpHaJ
lv/C/02wYki2Z0V6Xti77ih9BBzdxiW9u6JqC5JIPszsEG+rmzwkZmRUZkilU8Y38CgzfZaVzZ6x
+MUvWXUC3iCL+9arhztJJd43XKZm5iwR7cVX5oryj2eYw12ps2RxW4y6GlhNCt0BYPeYeYY1F6BO
k44YwzQSxK4fAEaiT0vPup/0Ry1B08Yfgdp8n3bldI+Wcrl1cgO/SYuuIG8DwD01RGXolhdF4RgW
RYdm6vZJ6zEIfTMplO25gyC3nW+ffM6fisXMTAFkyUDqtQt0+ASHBrSIRmrg2LWg9tfBRxUiI7j1
g/4zpr8jyt5y/g2jrNgS7cm4Op+Ddyk8lnt5B0Da2CJfk2Luc61uBvDfpVu5wuuYhnglMx3V4PAz
J0QUzyhMXtGd1fJ7alF8nk82MNR3AeEih/NtHrGpKCx0WY9HGoJMuAbHdBqouLvVY1c4yx7VeJzx
XwUb7JoElOAN+LaTA9u+SHSYtyD9IO1eujB+azxLO0AMQJ66xsjSRGFUIcsJXlonHiE94RhOovVB
ioXbPu9qf0Y0QENSEWfir31SpbGHlgBZpFx706q0Iw4XWi+8JMyjwI2P0GnreMWuYI/s35ENBtDe
ubCE91aVDUpSiJqPrsfz9WdWUqbmdBDkBIuKzhLyTALq9W4zsIUQW88+zHDnkp9lt5S6TEyFh+hL
y+BwteBrPtUOC3RhRTQBc56hKaXAQaB3VrZRwXsl2ELRzL8EXcUczeVSmwp7LcItPtYh9BAS+BWt
tk4FRC0cHHlm/bWOU0f+PYsAWf26DQ3eOZOw5syXYUeTuWyp48hmtjVBvzmy5a4QKnuxZU+aFH/T
Zigws/O7FmS0M3jW6w6eWQ9sZtGqRxmuB6ioxlpPvZu5i/YB3bJ8pyooFBPT0Q83yu73OpsU1IIP
5tj/fOADGZVK53FdiCu1ikisykKu0zcAwMJyrFveHIJUzOYC8fJrba42R/XHC0UeaBVYqSvub8P+
Z96+JMAfBwIXFPz0fzMBtB3XVb8CBPoxwStmh81TcanUwQxXDLKNzS23qwVOjI+DAN1L5T/+y6A/
GO/yfqGDbDzcswFGcdDggYArHAnpeY0qeOkukBprFjjJbukE7Bcf3UJCLNuLASoKuqQtwmal3See
QlsA3tESGeds05IEgpgjqARNYtFUmp/lg4B91CYS4gS4DtMUYW319fWSHi0Ixxuk/TEJvEaMSEJC
TQF68EfnL+NoW80d6fXgOqfrXKx9ZpehYa5IP5312Th4dcydEQZfH/ENIkTQUv6q7YAmMlhuc+V1
q8x8wQJZUuqBpAoQAHNcy6xmoNrpw5/O8ZgRNH6bI8EpzSAlZurPOgmFgY6Zmx/ZteN4giYiLoP9
yyCMX4tl2Fzx3W2KxkgHF9Snhzvs3qSulzwIFYJ4qizKoQ56AIy9N300EwPRuRV/MMF+VhdDjS9p
iE2EPgOUtBZAWyP/UNmmDDLEZ0IEBxxFMefTvU1sKS9KFCQm64yHHWoG2PApIZuN0imAlWReazQP
YfBbkj/0ehpgCmCeiVCrsTGQhTLrAdK2Ub41XpIakMiF15SvdqnkgOATJotDmTMcpHywFDFSQ+BM
Q5de9cvy5cphSdQGZlSNXP0+kT7q2coTEuAqTIw5DEVO+4GcaVsXQINyCwwrIpFl8x+CBYMhmgce
SwZuwG/EbfGiHIfUqCtHRbj2BVgYS9ByQzqK7GkTOkd5TjiE2iA9qEoF5g7MbQ2gRlSGilI67/nk
Yx9h0F4JoJ8fvwXrwFNkatX50/OiINhB7HSGrpQon2oSVgGMYGZMi0w8HcPinIcYxuJLBuIhHS7T
1EPZLkwTKz5GO8Vts9Of/Z3hXxb4AsBmcQAd5mG91YqVWnzGUL62peb45q6sI6hcfNuT/zmWCsuy
9X3VSef0BblorVB3KdzoAV1ycgFQJxDMGg8RIQw48FmraFEaRHGNBtAqQZSVbz9fCiGeFzGRx0qy
SHiMSDvgTePSExIbNT2VNUAQbcOPW+1Qrb/EvOmcz7oZ7arGD54BRTqdjsIqQsyhhzw150sBejya
bAmKT4Q8BaEYTXEygkzbsKah4VViqm7yFo071eJ0zMH9wknqoQoSZ1H2j3wKlyKiqd4mi187KXPx
2VV+/UvuyahIouxwSFj4FpZPFbrbLWiRwyZJmQglKZ0peKO+qxHwYBJjFmTVnyI/rE4VZXejRB7k
Lp/CocSaOuttLYY5myZcKXiZjzYYrd3c15ZtCQ/UW6mDq54TmXrz6HgzZoG5KR9E602nsIXf3CM/
Wncok6+9xxgW6HMrLJvdc0o4Twf+DUxpo2PbkJR/CGWopkrLY46VCGeW1+m2OoBjIIOzU7IwH+4p
rFYcEZtuSDtIneeH8Yk2Sh8KzLXAIGj1m2tLe+zQBwch6TXWp1yOfi18Z+jdSsg5rdw3l3vl9tnU
D4vyUjMtcGouUPwQ/oddyw7AW2NHvlxdZoThNV1VdfoMwQDc1J7rWPaa5naUS+Eilr8SXvqDjed/
lR2bpFT7WmfIsYP1WIZExDuUt6/4zfryYur9eTD+xmaWm8BttlrNUwTUtqE0mfyMdgk2cmNyIuLM
lsR/E3iGtucHoBtsBO0VFO7oiGmem+kRNZ2BSoRVc7l3vu8WouEheDde79nFjzQZpNm5Nnt5oURs
2mCxlR9C8M6hY74IhnVJ6db/D+Dy/CR9toe6aBZEG6Vm0KahaBQ2F6LFcr9aFksWC3wYb7kEs2/O
N0BMbAZVO+TxPbPOms0yKA8V5TbCih+vKTwpdgGMFPWdDMOIGOncgl7g/SrUcJfTNItX1I5siI3A
tPLkFKf8C/unkwgv+njAzUlaI1b5FwriU7Cm2stGNS5YK5DAGKQlhEH1vkEopBQKxuOWnMbV91gh
pyUy7ani31rznDxEL77sr9UhtCdvR2EEFgnXQ9rIzkpO3lt2wjcK5mlUZxc+10hfd0tl2+J1dMzu
WPyuEJv6NWNfd9J3KqBK7BHb+wi+TQkJXS4hfBFn/jiZ6YZakpp/gQXyu46vXOpPGDw6uAaflA5/
DlfPCpvz2GjPiuBYqqYGf9eRoiQnjymfd4XaW8RfyTeMwKmpzqKn7Z3X3PVtSGDWSlhcJnM1vgLV
Xn1sVpcX9iaNNGf80y76nQplEvMtITQWPVTmgHhBdGPQvh+zaNhhYTT5bHu3lnGq7O+ImpmQG2q+
/8hPj9f5sBiIok6PIAjeigIzMYvEgSm9dREjUtFgzPQq4aKyHkY0dCKC6bCEk8FmVVF2rc7mpoGx
Hw+BMGVRh8gPkVHVVY3fGg+UWPur2jDd7s73FTB21DQuYiwTLn7HYG4YJQQlE0G6zz+XK2Izr+Pq
m7kXCbThc+uhmGsKQS62onV3jqSjJZiNN3q4JII82PbG5yUzubJGWTcnSpTOovC/JNxiLO/Qcwn9
Td8eSkzDP8/imZO9pvH4VUUfTJtBDkKhsCUWCbPhXAc6A6ESCWgPWKGZ7AudI2bC1hymYguk1eiK
sq6LMguf5gMwv8GiWjhS8sMyN1PQYz/FsXGytparSRIPv6xkxvaEZV5Sjsgzp12NXqXcaLjpuuWP
zpKU7Ic9N/CteWZ+3RiQk6PpKB+FA3kv09B2dkEsxAVa45HEO4jVJSBauIJKQTIpRYdxnIOZ47Sa
U5f1kojQBbS3ofQPKX9fWvygoNaDSMk4u/iqelvey8M08kCfuhIH1D+v7NW8JUf0Bg2yfU9YbBVK
X1qoXQH0DbStdn+zvw8dOOSJ0n3HKfN+blI/KCLF5wWkQJqzweZ7k7mtEQz5rtujtfpbzL6nJX6v
DBSFBMdeAHcCStz3q2cvhKwvcvw2Dqmj955ulvUXRH8xaUQ9FNZF2TBaRrK0XGkd8SbatfGHc2TT
589dADuArTol5YRWiN0/06JTXwqbn2QJTu/vHJY3TXbqq0JGSgh5I98ZunskOhzUk2oo1hToWUYY
lFi+Iunqtb08RF7dwvxZkpEwUMYlWh53zWsSo1noA06SOZhleP4wBmET1DRCN2YPX+BGHVZuaabB
MUX3lWlTIJEDaGgkaIzouCnFIl+HvNOnVU7AKsD5R2cLQiGu9C+XykfIlwPeCtYs96+1L+sow7k6
JMR16ZZDqDx7h1q7YkU9lLgG8gaWz1k9SE0aVoldqosPaZo7lyNl6Wd6mya89/15p49oRr4qKxZF
o9vzMTL3ubuc8D/NCvaxHydH/ZidVxPA8W2foWQRHXYgpwD2VFo2m9USlUpbyDzwDooDypn/Y5ec
NKbGtRqY/eaN2VU8FmoS2ez4OAPiQyvJHfS/U8wZwyqtj1yZvYNknLUPu0XLibZiPuVCyLBo72DZ
+oIx3WKjt+kTNT1kfUiyqBvTvmdA5niTxQINDQvjvZ/4BqlmzhQcxsKidZxSePxYnFB42xZ5pDFw
IEFl7GcKIQxBF+Ekz5dGcyQo6RSOGP5E/oPKvjP+/Rfw8RQDBKEO3pODuqdfOrCe64NmmXIE4al1
5DiStbTt25bckbIqCI4+doFdnJ89NYmhCsfZMXqDEDo43XSpGAw3LiGCSpgEmVO/KvWH8+KaCEfi
jCXgocYb1c+EktW5NTeo7qj/FDgWy8ConOCwQN5mvUFZFXbHSavTlatGemSigLaxpvMKwkLMnsCH
r6pwlHVEtMYhcaZfnmaAR2FJPsNV5CGXgtPEBY3vF7g2Sp5BFMXdS9P3gkysf3HnAVvj30hkRh4u
zk2ahzoTvrWUfrZZn8z9j8/AQlem5Yp4vG2nQAbNs/ejxS7NbGFatmo+K4USAcfClyARpSdu5j3k
/F9fLFgeoH3cdbWanApMadEdRifoObzyboU8eplstl17dJDbVx98Rul5ZoS1X97j1xv1QwAP8+JG
RyM5AQVjPW7k676VDgqlDdKaVFK9wpEL8Xs5ElUwhIaEnTz+ZVtn0AxnhG5Z29h9sD9f69ShRC8a
9Yk8CXhePUqbHYBTB7Suq63cr1czLgv0NkhRpQXisz+vGLXZILL/7fsaCmZ4a6nJbJjJyO6FrYJj
6Vh46Yk5wRaiDC2ra7UawzvqbqmpGI4c0bD8GYr9WFBWfDkXUvCoIemUeB5Ki6+ovxj4RMqYXfZj
9luZYYwhtGUpdKzCwj0cyLin/sQC8ehYI/CuUQlZMBvNhDa5LEIoLf0edK87nDwfKhBI0zQMdI5s
gRMtUYf5akYfWN7CYZZ8VVXBGxuiTcNfCzUqcZdvzYvdW+3qDHtPZHzqRZXjSTBkOT0c5iDbLEnH
5VGVcUv3pdugtR8hEq7Qj2oYGm6yE09uZVA8CEWZYMAWXFDn3Buynf+tspjyBb9tB+vpDDFejVA3
jDPVQKbLiXjppTpfRxKUdbxCaE8bICG+9IOfbwYp5Ym82oXGDZ5YN9VoCiRqKSs+s1b8147wM4Vx
OPuhITcEFyR9H+96BVxiLyQAMzSbToaPr9zHCFyLhlQ0Jo3WfuosLz8gN0Uwn4fWGaCQqdTmmpLU
aiwGswnN2KmYUz/6PAxEgXgpmmjAQiMXMrw9cxqSqQNdS3EPHYICEkZ8A5jvsZL+rRr8h617yhID
X8W/o7T2TAsniVYu/GahNpxpSbs5XRAEvg3FcXsAzSvkAD5rlkS6JvKIeoYsyMxMOZjEcpyJFayy
4KiMv9xtGwEXNkj5WvDM71F1ubCjipPVVScrqhl/UmJxj5eNd7495qp/IN+jkkXQtiWop6fb2Cd2
JO5LA/FbNAUb9FsU+fZahXLmlC+HiIUrieEQdqGMSbrdHIrMa08CbX3QTAiQFoRWTXpSuoP7SlJh
izAysVQVycvIv6I+a9iF0ZJtDB8XHQ83NNCrk/c7S+0e0Q+meAAaos8wH0Hix4y7fQOvO443bTnw
kcYVIE4R9sXn/awEnpAXq1LOuNPRMU+MkVKwQzsWrplNa4nRMplWfpdCNDqKHweMyBTndpShQ9/p
r6jzEdc0MxhWXCb+AGiK8wt469d1BGP94vMwDVO4Xh/WQhTKffPL55noJBGC72RWXyBwSy/vwb7E
hYQtRbgfLSmQc3Nk69vcWThoI1pV8X4jHnPa8MN7cTsK6VRMCkmm6JfILVuaBRD+1As7yv+2YlQp
5yBNDvLI81/uxcltHiF8WTekQdFxXTcD9zzFHrlvtiBo6+4tmt+jkzaoZJ9WViGKDZQF5Q2ptz/y
8phv13WFcXsPKkyW9BJWkSnJOyKjZOtlMXIAj8ZjQWpimYbdLUoubs5RO0NttsgDgTQkR7vEcT59
bCJvZFkFPkDH8quYfozzZMH/75HJkq27ksJcgI8Lw1XD61Rb7pzxIIrrlJDfdUXIwqzrzZ3dFJEW
0gDevLidBJ4MCegT8nMuBAlNRn2KuWKJd2HDWVBRECqQYHAudIyiGbJU/AEX3sIpP6c1iQk68gVl
92xzIdAhp+iuh2e+OVRmrnYQsrdsdxw4hAxoA38mjPhWxl6ny0XiVEzXwHgT/F0Lvat4GikgYJZH
zRjsqtXeuqCZOnxlriW/7AWIua0FY3V2U/90pXanWW9AbT07o/9uHpC+KcJMYXKD2n6ZxvnJJG2V
aVwVFZT/W5AJK1QVuhqs80ryyRSvtJbkxW68XbqRvycSiGW5lLnv+IxX7b+K577+6pi7Bz5DbtGp
7QXQqqD0D8LVMO5tx9yBI0Z2Fg0oacqGBXQbLjZwDzJJnYlWqCgCiEsN5ogj5B0dqKnmpobvgtOE
HAg1kufYZA1xFmnmNVijbJuXCVCvbyIoplaPfIGu3Ba2+SLWQwTmAak7QQGsg7zruBE7GIyzHvfb
6v91LAzvCtwE9eafDPcNd3RV+tL9ohGpsMKot0AjeryokRPfhBUQEpJeC81kHxhomrRup38qXUC1
ymi8x7WTkUfFIR9VSLo5VXs++gRk2Xxyjo4Ol3MV5xuXvX1ThBt+SmO9cCIlmnr2rdn9qYKVDgws
gEU12HaQpGYpUUazVPHGJpFOylcj7QJV7bjnKfTfAcJKxaQMS51vbRtxp9PLNPs2/v3FIQgtgx2Y
s21PuUcgAqI2JLwLQw2AY5s4cT2VnzvMxUE5hnSCHkA49+iFT34v54XCrzhDxKERTjYqxL18CD/t
x9acTnIaVcUYbVCtoinO+mQzihnoa6Gt7Pwjt6RD1+gOUwmlh214sRaUSzWmPtuPOr8GOw0vxI1k
VgavH2BmqL2fxmwo4SKpi8Xzi3tPjpKbKLCo4NHWkysY/gj+7mHe1zL/cRSs0FbYHpyOVnLf7Kye
8TZ+KrVgO3j9af/QIqTP9YIomDB+w1hRlCVxa6WHOtpZ+ptGXSsF+dTBjhsMTahz6onuLQfsODP+
2Dv/llxv/5a87kMvWQF/5AA/swFam9pliV44lss3bbCuuFYLrHjrSyQ/2xmbrbF8qcfQl+Rf+O7M
AIwy6xMqQGp/exEU3GdDqpns5lK5DfA0iskH3dpCAstAdQ9MrfDmMJeKem26N+XgpXm7mqIdMLGs
sPkNHYvJaSoB3srfDVSTDAhL8yaTr/SIt6hxpIzeYgk5mdrVvWxatutJ2+n0etfAIKgpKW6AviLd
J3MI5hZuk1vipou/afqVrr2t9fLg7VjxVJI6c7CndWMqal7KhGso7UoIM37pfsMyQgwzqreKwDBP
aX6UWDY+yfcvbHuGqkL2++2uvKY04/eXDv7riwYYLYJ48h0ZCHw8+MId4qH0z31wPRplW/ZRetti
djbL+g3sqXwP+j+ir0ZHi8zYPiOAHJESU6d+6897I+42VpuP0PuHfF4nroq2vKdDxO053Pb1JvH4
h3wgX09tw9sqLC/cxvZVUREBya7EChtFuIJbtdM3xoA0i0TFLfCg8smwl2I3lvn/UK45vDOv0s3x
lzz/7mP1H6vKJhiiziFLBFM5fzc/BgSX8gVZ0nxc1pDFq4TjTqK8Yjcc/H9uxokhJbkj3tAvxLSE
Awi3TBZpIc14N1aP3Fu4+h/5/hGMpquj19WGFERUPobZ2J4HZYq/UDwj/TKFQ0ZA3L/xtgjEXO4/
3PvRe+HizbD1UILK8G/gfgiQICWBjy8EsPgSRXBu7xBkUoHEC35zCO8O5H/WwB/Xt1vWwWy9Q01X
xaugpLFaXK0ZWrQKmlOVwjwvKwf95bC3yGuC96A6+TLZmVUgUwHyrLwnkzs9+eNyZpxXtsNdF+Bn
rZPVgvk4Zl7Oy9fHqtFBsl2EZUncjoWuvf9PL3n27wsnW2hofaBGWsXyB6WsY5TJ6sQFLHBKbHy3
ch7lAP08dWhadyy1VeUV8bhX3u+Bi997YwDHkJnF5aLdIV4SxFiz7YI5hQsJYQ58QfI3uCv9D+gp
bN54gda6oTOjCsrD9ir59GV9TrOnC7yrpT3VYcAd8F2+fweTGfp9fdjAHWMC22RAQ1x1c4WzP9gY
ZsdMoAXBGOGVXCF/0LdDdXjisMp8/5KtAG3vFoWlP7Nn4UrEPwYLJMS7esZ+c9RITZdpmoBJePOb
PIHM4VI6mivDU/B2sCnqRZGxSefr2MEdI8IKFQGYVMhTAUDHIF/jeAPybWrosQ3wEmXh2GAtrCVz
L9USH/59c6xHha9iU95/+/OKauiinmkx5NnT/rYVg+uyi/vIb9kcdgOK8lsLjVUvIax+l3pcT9V7
Gk0BNnpVJz0r+tUV1ivdGUGlP4jUqnU0MkAvpQ6RUe4/nm2lCQRKdf7jvwWYel992PqhuYPaFe5m
DeGPkx0+1l730nSfntT4oKnUD+2RQRXBSqqPvsRneNz39Wl2FoeUrSroMnTQAPjKpKCMyN30X+Ta
1FJ5Aum4N3me2lPW5oJP4xbg8FMkGSFTGrkSbZwQEcCCX3KcEzPH51kVGg66Lx07XuthUkWHV1QJ
PqAhos9LNe06+P+KIsyUDECPHKQwukGRaoF7AkpQZ7g70raxlvhMBdSX4lLHdIw2yOv/QTs39hsa
nCl5YFUvD7+E7mu+/c4gPAIFBL6dXWXOGcrS+3m+S2FrO5LaolycCidfz9COU7hyx2gmOfLx5PN3
jJk7UxoWp5JRr8uMPxFV38j5c7SRo9bYogMdcPvFVBzbBdppXsufIJfVDDISlaYTGNWaSF+Zf23I
4fy2Gqpu7s/3NLX0+1qK2p47mqHFQ1kTdGBKE4Zd391wwNxynJ0II9XWFsS7N4k3GuVxPpcnI0Iq
rChy5u6lidvp0U2F0ojCjbQRZDi3roVEs0Ud34Ez7TBAetS8ZI2YbFhzVXohry3wfggsxcqBc1pG
GPBsw8EueFrXLO/5oSXg+htXOapEV2rA9Bu7Kdid4yiTrXAQE9jUNf8904ESEjaCSzTYlyO1U+uw
jB8o5n6MXVqf+nQYe9DHE9G0zUzP3Jsib3UMto2AEVrhI+n6/cjtFEEVYiSoku5xUDnBIaQ/Ps5h
7LfP8o+MXnp8syvJTQN6aTgP4MkQuTwEbuwZg++eqYbyu+3w1kjqlT+y7Ikfzk21Ofqfs3W9k07M
RPiikENamilbqUngXHLuWilHE6g9S8Y/dW2OO7egRd6a2060BQT4Ioh66yJxY9vjvC7uVHA7WLIw
Sa1OrjaxrrFGh80x5lOToWGuUsOPXJApFWRHn0wHROxqimYb2JGPz9Hif//8xHMMvGk5vi3mdTEN
Bc/k2bRZJzXDa3YlDn0MENjD/RQM4MOcS7dhGJFnyQ0BKHO2K06ZLh4beAzsdQFytKyM3mug4Kx3
ZWHZ4emIcOWvMsDcddZ/tmezVeX+IbNJ3Yl13ATF6ScQ8+rC3Mc4P/ornT8qxph+NYjKFn8c58Ac
F3EaG2y6ctWwjjA4+iGYCDRrYhdKd5FzawzlLqSR2LtCy32j0dvIAovCw5FBskVTyfUx/zfZwXiC
6JTEHQoDwy6w6FHdQF6a3+UuXszEBAYNXE5UpjUrU1/TZePvgFDtXUqNO51p517MwL4kP1W8ESa9
RUnHha59L+IwtJE7gpG8/tuDEl8KBdD2PBs1HWvC4futmX9q5IEzLGGbWEOS5r2+R5zAT6l0jfCb
vRhJFzmHyHZ04Und1SNssypZxGpympr/QYo1Cy3GsAEVXy1p/mEOS3zXXwPusAWg26im3n9ysHsQ
HeQY9bqvPFTphYa0Qwag3sKGCQajs92kx+32Am3a2YqaDYBZtCraqTlM+O7xej6sxoUOuBETtUik
wtABXvVqvyOTaRXjzBKxCI0VryKyugJNU6zrxxpvA75XUqWMMkyk8MS1sLoV7lBAqkFTlN3PUQNj
p4VaMZq8p4lhhVSS7eEkasBp52CeGaC8B0qx0Lhtv5f7M0Zz/Q9k879duWyoKtU+Bf6as4Fjdizb
9WsPfgWD2GrZW4WSvDYcsMqp6514nQv208zEAVv20TJ3VCPPCgkJ5pmr2bLBnBNm4umvA9pa+sHV
c1+GbaxsFXkDa0uVPyW5cw0i/YitYGFYdqF4FLmoP3LwHTMU4qjqfQlQdaXfbBOK8vaCQdaqT05f
aK9xOTm2eI4/ENQR3hcRxtUH+zzpMKtFZq9TtlI0FR8dpafDdA2gyUmT19ogtiwqzcOuP9ODWPF5
jVtWCwa/6r67Fobk4XapJmn4xCodzdww75SZIHv4AeckZfbgIT78T0Xz425tDRAYSdfsKkSIy5nB
hUDoP3nZYjVEEBnamBy4kGs77DhCnvzyhwcyYrWhbjpElxZKbPo5sz7te6rco9AEHoYdTNWTa0ql
FtFJxq+Il7uY5AFV9zWlN8mc+2NfunHJ09RcXYAljxEVLiAf1MeCH9JwPE+TwNAouUyulTWFClb0
Tnclm7JO9fSJQZAbhmlHea4P7ZyaCjA9muN3wnSVIK8IR6XIdGdYXYO/vX6uCEZBDd9wYaFBN4lq
7jLuz8bGmrajkdtVVDdHr3E1YPU1A4DQKSD5IkOxwjO39U3NDkm1+KCKBZDH7hHmMIXz1vlBS8Hp
zrn1SzZLSXzA0fgR1pbTZSbmnDpSyxM1SIQP3rGRhH5qUilLkhczEElgkodvh/YpCGBc8SAALSOS
cJ6Fkp10YaF/B+gIVA263Dkc6OguetjrBhpCTrX+aUXIn1H8gkxXrAo5o29+2UcblbNCDzcwOvLA
lTgv9eE44jGXiqG65MTNKFrOQ7mQZa+GbBNyucZDRe3dE/nMNgHSDd7AfyxDhIMOiQFWTmo/et0m
ytWJjAIg09uCK79yz8v7tZ3Cmdi/CZ24n2LtUxp0T+eT5FUDzEtQ7eafOT189ntYbuLqiEKquLOr
BGE70Sa2cd2FgyMBcreRZA7H0b2QLgAU24YGxmRk6tQOrPogt5mnOLF8TQV4VQ4rzB0jYNem8e32
RblpLt+qj9D/NDOJ+A6cFNDMG+xrCFR0bUQU3qQahQ3xF6MkcLtmrX4yfgnMUJJlONtP/CV59kQm
1RUdwA3gu2C3+7e+RM+t5MxWDVXWyCMcS3IJwbG8jO88Ej6WedRnXTzL/2NclML8W9TQEG3EnnLS
SEAXlcAJ9uQxF0+W5QzpNOEI8uaxeXxLlhwhLJP/ClOwvsllFEO/qMBqblvqbIsuZd8LunVgkYFB
ashjzdv67AIj+yTswKH0dkLecBSp7M9ihVOPqzyJJsuTk7dHqIyPqJ9ZGm1uQzpl3l385N2u9Tuk
l8bi0omME4XSnijlb5VrN7YjLd7eu6b092qiofs/aZHmUmeU4tEG6utjNtZmALDBHEOoKOdhA66e
JGXErcWt0lbVsypcvTKzgg9nvio1QT8mKgmWw07j6WfewuHzEv1InwcKq+blB1McupFWlh3BDrGV
aBsednvXfGFAvnhtK7NRxmrpOAOlDm/XtuGcv9TTwx+U3E7fa+Uisa8iDZbSA+dUbAe0lxZYQNC0
A55aC8+MsKInNXAf3Jfz7SRUhpid2FBq6igGnaAc0JS/MKA5G6yUwi44+0BBkg/C8lUhze5pX5fn
aBOq0Cfnj357RcpuMwJiZTAwmaW3RrgrB2ycAIkap1pwK7ZOMdNWfmb3o3e9CxcJK3xUwC1bGwL+
x7ZlV4soeb5Xf1OUa0iYjz4wLnzNavA+KaPrUCI8TPSjxOcvkuHfdL2sbkqkKxtkFWCEYzk/rRBg
2A/4ov+EMiyx8/pZgDmxsSFcmUVQmbmDwO3xOTJNbP1InUKefEZ/61sqp+DnPKKjAAhftuG+E+V0
oiDt/zRldFdY/eLvk7dWYIpLOZjEd6IKWuMn/Efi6SQw1KVYhVQkcs1tCBoIiASDzmuTeBQRLS7K
tfdKa2Vp3WVQ6i4EC53dZZyHZY9yLj4ZpFNY70CpKosJ0yOGCRXLyAkK4IeTdTjFDfROXLLiNojV
K+8eRDAmj+uIFdp2LOgzVfvzGek4C8FRgvKjQbRLX/o0tYYUZrn2flMnpz1EoQH30CBK8ZPoh5b4
trUTaRRqu03eM3x5/1DEdAu2TG5094++xVk3hwbtNRMv0+hir9cuY6Co3ynSPCxfj1w1UEQdKNmA
2rMZQsRwMX3iepskS2jnJeYxlhf07OvRoW/HibL9ZEnvqFEtDZgAGXM1H1HjyZ72M3+ZUrXMUFjO
5Ofkm7OCB0q+lqWK4EtrHhshMbXmCbCtXYf22yrAZbyYYW6vRBOceNmzKQuoK61+5s8PSXVF5RCh
+Owd825JEKemg/ZdFNsvY+HKeM0rKHrxkvbx41AiZ85eLIhILWCBtpAINvn5c434EfoaMcK+++a4
O5GvKbUvQafdUfsNm3ONs4kr5PkHDafojsO60Qgrgm1Kpqe5XsxmKscqH/XOzq386ltayK2Bh4bK
/dRzJA83zamcpgGK0vR7WhaRFx7Wu8GM8UcXB2NCqJ7p9LGcgkoiOGxbd/0eOnN0L2zrWN4F2mmS
XRVClxXmVcL5EvdhElaD63uD2gpfUUHXIS93aZF92smGSi7O1yLB6+nStB8RsroFFs0ZaukQby5K
bOVfGDqywc8htnszJuULrqxkw2JduzNVfAu7+kqXUezjUTr4UpfPXHYUSpqeOw028+sqdb+iirIu
d84J2R8M8sA7lEnRjiRc9Bj8MQ0TbT04cPWBXeKwXB9c4Q/iAaKwqmTbgn/1nZETf4mo7Rwop+dX
hAhKIbdygjH3+AsmjhUp3jKEI05PO42IV+52R+wQ0SVVZyDbj3CilT5kRjNlOgKInWvb4lQH8zGL
e5ccqcWkm9xO2T3+dw2ilXX7jVX+GPoXkNpQNMpLDjxPd6GHLtYMXq/Ps6KJ1KdouZxnlMwGDgiP
D2L09hAZMWhLIDJeQsVJgrugMJ2W7zsn7/fWV/XkWCYj+C0UTPaVQ7KawpOXu7DRkiXHqebCDht6
zVtZHgbKxHXfzmXSCXaIvpWOIj7WxXwFGR4ulIen23sMzYh04lCr+9JgatGPJZzpgLdDi+qg37iT
vnsLGmA49Aosbb8dHtYfQtiYMov/aTUQsYAIriZF5HKsqzE3BmnjbVhn2pfnJ2Xbji49Fy/aw9yc
PqwzpEPqU4MgNUIxYUAeHpDDaqIkf4LbOd1F5/+/CvXzK7FUxtyStql9l9OhqNlFdMC6MACFe8tN
JtBBvFwba+r0jON+apxKmUuvFN/9NWYuGcmMSm51ycQnzIdH8Hcgv4e1Bt2ENQTS05h6aCl0huE0
Xs60LAGQB+3nUJV7SvPYI0cnxw51xYkJoX2SEyDUbGgvox25KCbMNI18otMMcT893s48oiWaZIYP
56kkrgHZYSDHJic7sj6D0V/jG0fTEQyIPtfYH9rEHXdFx0oaofoWSuB7viQYCe1aL8A1fozh1qBR
+GiOHdoH2xmH0eA1QHF7mzYhGP3LE3J/aTNnVNy1IGiZWXzhiZk8qwlwniqCFzb2h6e+DVonTxBZ
EOPqvbIeh/Sr6SgSe+1+BfUX3GjQuEIk/lkUhMe2ps4Ihh/hPvrZsHvR0saPkjC80OxJTmRS9xPo
9fqqEcd1ZGXa630Ot4APzfZz/qrE4z/nZK4wHo876jM9/5yvkppo+KeNJ/dEXzHU60wqN9kRpPnW
/waQj6sqq7+O7jvlgzERzn9Qus84YToXOmLjiud3RCHFEYeWL/p8uwGUJ7adUkSS2AaIP0lTKd5f
DAKPehcC+zkdnoKZlPTD5hcQNTrbLzKgsWfyETLjv/mvW2CZ4aqcz8Ut8gASrdZs/a4pADeurZw0
5P9BtPyGgg+f3521pRp2YphzhutRdVLCPUbJHY17Kw259XW0UGw16tq6lCnpA9Jd8Dw6zRyKRall
MwIXF8KOE2lMV5HrGmtk8REyevsTn+5zth9ZtwLkYjXDl5+8WLkUGr1/c2TJb6cEGJfSI9motT8x
DUfVZUhIpQuX+2NNgYx08sQSBqirt104/2aL26ykRder5yWLBpU6Yv4Lvj33abi4slQTc3mrPVEw
AuRgU+6ni8eE+YmaZ3hamqO3AWrMnH9lnSrVNvRL8GmKXXJH/d/cpU0NoS+1qbqqrqA6wURgRSzx
CII/+0S6aDGnX8Lhz3sDNyaAK1OFcgtPam71gU3at9jA0exe9+KjYKBdMpPsEIoq+Gy3HwtgFw35
9AZ5x0IZ8BAtfbtEiRMpHGxlRAF5uQbNFV19EG9ncHKIX0Ooso32gy3bapaufGWYIDKG3NTeTZ4N
R2qB9jVEWD8Er9XctDPIyyMVklPQuzoOBP00dWdx33WwmpU2h7pGB4FV3OPVYfBpdoYVkin8J09V
jv9RFueRnidlt/QHa0epKS5rYKhft14qI2JKrySgZrNbZECctHEE3Y3racG5twdCVMr6Lamlf2xB
AP3+C9C/hlvQ7qxEwoBTEFSLN9W7WYkN+mxkatNorI2CAtxBkqHnpMiyc7BCCH+A9JrqRqYGiJ9X
QWTq0f7LfBosHaA6OLOP2D09dmuSHBj2yJVSBhykaTJiOQPwTgRaGtJUiE2NpufJYFBZzFYVZ5ik
gmJfn5Jh4E4m44HMHmK6ugplzmXR8w+tk22mn4q0grAqXdOl9j+ZQTUUM0arCVvhaeb+kcErZhgC
4gsRuAw+qLYSk9f1y2yJ1H/AEw+46bXM9mFrX7K3DeLkyte1xnKFP+JFWY4eWsacAexqvMK46r8A
xmDzPuosn62Xs3H9Y+285kr0sAijUm+WZxy5Fo8YcO2d3TxP8VbIrOSEWAZLkxDaOJymvN321t+e
BKT1haBo6gX1oWPpuAD6+bRAIhRJUc6nn4pyIRsHoE0AOa4/YDjxmF6pFuVd3chaFcbaYQq5JbxZ
19B53vZ6BDFiVGp/TXXEunHLvX26cxhMT6iJY8q2n5wrSgQPJQcl97ISevtwyEriQMNT/DWrbZCf
DhheVdSyWYzAAO2i2wm0ByzGel3Whs4IRSGxU7LebinrLut2gJFHNGpin7zqq8oMIWWYl36VCVsO
fGtZw2iiu4tSe9FqPLM7kjAdJz5sc4Q1SQ+UfysUWwUIt+vEP4NBhSgz/ZFhUMx2IaV5LbzazRYq
hTHUy8thkfE5aAoQch9Bx8R5R3LKymrk2L0IMIHOgVVhJbmmVlSSigx4/fAFMIYxDGTMwxSgOpsY
URBgWQHQD18I6+iGypDa6U7bOwtfKQFWZm+YvEADIL8gJ8Iag+oDDufyIjgZdcwaWb7uo6PuiCQq
b+kgb4HsWQMYKFD6WJKfs0XX6pmF6zggfBA9J2H/WkqD4Y06Jk8/6rYkZK/HzZsOr0hSfcVezZGn
3sSPbfpcbU8fkFQ01+/pTHEWw+l+BnIyzxpRb5pB3mo6IMXgbCMH2fpPt0bAdABX46ZXY0eVUXnz
b8uczIfoRJqxRlpwcTxu9tdFS/KAP4zmY2NnAMmI5jIm8wgdKczGEjtGzh6TSWdFdZKDfdXJQ04f
bcY2CpJtiFMOCnJJprhtrJCkK8AQdabSgf6nuwZYAPNK1AOgyHqAc2r1C00hrKjgtwxZ60iyhemO
Cafbm887rtjMSeJLuqGSEkfsEVTWm2nR5ENIlPoDiRZx9XxVPMhfAWasn8ZEYBkQK1lvEjaTwEf3
Dg5bRty4w/KZfUmQuhva/SEoZmvUoXYBt0DQ4vkrYUAyGMsb5t0mGhOBj6lkolKLO9HwqhJQ1hrj
tKI+vJn1zZ4G9hZIqJT+oNso3Od2hCMq5oqLXaMMFoVcym+WEqd6uZ+noAevQXbOZTYt9Zj8CCVv
e3c24btrUoshiEXwzesQiA9yxEVfJw8v8Q0wOsqw1EHdtOyikNmrtYqce53aT6ddMpzX60Fh6yUG
Omni9AwWw+QcM9I3qlIqHBMCHmG923AGQS2N71AVJ83Y6Z7y4C5TVQjcRogQl6KKTtasY/BsHMCH
mpx0dqo4AdT+bDPFgAX18hsc9+DPVa2w1Nxd3upbuF+uK1U18VuTdsYjJh47c57jYxNpsvFO/+hP
hxhVqr+HQdZvTmh4MUGSfSiKNN1DDxEZfvApx2iFv+ZVWBzoAHc274WttNgia/AulFk6HhzFJnwF
dDgiVmiNFxcnZM77b53BDBb1mk3dTkFc68pFrXlbR3lk1oTJ80dnC6pPgN2TqFpLTL6ElPjgJnRP
0J94dNIt1GAf4idG3QPmfNqznbGeVk5FNIl6IlE6EPwXvwydksJ/ZfPHf7dA/aFbP5tJ7iWyKzWn
d95tCEqfI19FkN8h9cp6vzeu8j3KULClHPP76+CyPLYjQGwBr6NzDLHupl3n6+fCpgFUb/3nxjVt
RKXBNUUGQ5ug6swuaySK7KfwNbdjuKHoY+umQH49XIPi/0k48LSOb1e7Kjb+AOYjxsAHCA7/sFML
13p7u8zDC9wRd7aHzTZO2xUvXJ0eIm18hejm3Evp2nwLyLUkPeVe5qJVTtjNIj74WxqWauMURCcf
WNbSTUIliXlKji/Hf2SNkeyIgtRdeqDy3TBp9sNcZ11uYYmg6mca4gpKBBZIffgycDsuQZ2fmatJ
M6Ar225elJgPG/d9YllLZlH7o12cCUUWmGGcpeGM0DR/a6hBKkmuUtLttOunWfHGyaFiSoWXOvSH
F6AUVuUojqHFcVEOW53z+p3rzf2ukk9i6NIDb6QWzwZxKEkX+i96pEM6Q0iZ3Nqe6WAIOnTTe+91
cn0w2WfRV4WCFIj9A6U4murUhNnu2Ea5qvrPVnBPLQdpTElWmCkYNIDUcIucbpDpzAmDM52aR8BF
414oHhZHaYz840dagvdo0ceNkf6hXo8d+78MMjUrNQsJe+LSfR8ClmQOpDLXDpLftQ6caBg4Abzj
nIoKUOmQx+ywCujutwfMbHnLkQZLPcjC7WTV2Oj7PqoYpZNqVOcorrxbLrP9OyYomWqabqw4ZEmJ
fiu17ayVRX3DunwK31/Sw9iDWMAqCT4Tw3FvWooZuGrdlMzcTJlLzgAPjSYdsmMmFj0A/odGDPYQ
4l5HBbnfJ8qEwkkgS3Lrw60+2tXl2doH2wD3UtqLi5x7y+Wxfnf2TH9xDtnG0HmMjyMVUKYVYGrX
B8kNsxG6yJ+z2fEbYeHc5xaZKLjdkyDVGo8QIsU7cmQbi5+Hg67P7kbMnLXcjfapkaS6ys/4cOQ9
xQk658Qw3gEoJq0ewd3cvd9IbIhQF7NAANnLM/j54zpkrV9z+DA4LwpzcO7Q4bUOuOgPPjjt1h9/
zVkEMfDyJVm2HDLzfeL5xanqfxr37HZWITf9xddhqP0xK7YAQo9LK3ODXMKWSLpU7CS5+GKRg5iX
11uSRKJGEpt5waini1q4Td55TOYh1PYnRhKlx1OJTzlitaDfZZ4ZzhvVkusIUQ7Qu+7ysbi/tcuc
sgpfhC+sJ5TstdBS2Ijfc+OB68jaesLt3873Js2gM11lJKpAWVzeJ8JOhRaE7PrrDmksgfI3h3n1
32zZzVXzhnkXpHz6HkWRWkLjFH8Z5oXCPRY4aLoXgSzj7g1HFQ3XK1Sbntpa802BriCyXxzVnXVn
kg2PIlNFvV46j3/zF4W47vikMNGkucHdUTVlibTmTSEpvungZLFJCFr86BrvMxqxXKiqqPM7Z0pg
8GfF90hZJ/3ebPQ/AQ15GgWCfuto9caJkFKYndqHAqyNtimmKXVhEFrQ2NrHfvi+pF+kYYuNDRhh
h7NoSA4LK7S9kTMSE0Yj7SI78bcyixrPzB8pOeCFu8Ddw8Cm2tsdJ0GnNxZUVb8zElbrdHTjADDR
NnrRU7WMX4r2sfgvZKc0LqLHIuG2P3UqcsbH0jA7AKzso11AbQLzUvolEOq//oscacDcP4I0vLER
7ZaI78wedmbcfIJjcE+A2VhuNonR+qI6XeTtBCkOCio0T8+0ShSlBRHi6PHDndIkWhfDQElLzxQW
btDynumLFRCJPllCGHk1bRj4sKoKmG+O3ZT2PLBjGCdTAQwpAJ/OhOdXm8Zych5HlCByW+LmbNOb
gZABLEG4LASS0FebqZkO390wN3izE48f+Zza1KVOuBW3lUJajRGcV8iZKjzadHfaCSkMn+wywsX4
AMHdKmY1YRfEZVxWAPP5p5QICedSVhi6jQFhEKNF+k4V/JkHuRjT8b0q2c8zmEpiuopnqVzge+k9
f9ITTdha+7laNZFB8al5j0YruQiThniqdkOxsRhWxSrsFcJKX0ccChl479U87/dt+bvw9wtITGJO
z8BZ95D0k5KpZrGdG6nUb1ofN5s825DoREAgQJy8yVkeOHGGdJ0HZTykkV9kNkP9BVBHFT5WTrHM
8KejiHqtQdqf4dkoUu9KdvJZhzQLi8KxayPkAE5CrWZKPLQPXn33XAjQhOCKyJ8XXflEUaid0pVd
fh+m56ngFcnB6Q2OzMQ6VS6MUp03OlUJKGOKgCqbRKIPzt2L0huGkkZTDHLGc3hx08FArgMR+z9E
r7/XD3ICJqgzbewwJ7NlhQEFLXYfoNUHagHQ91WAd6zeEL2/52Wz+c5DH8UJgUynHxPrAm3huwa/
fzgxA337c33pU9c072nB3W6jg0b92uQX3KN6r2XzoAA5pbd6B7jgxeCt6krFPIhQdyhAUd/FFLob
k3RWbU4HTEqdf/Q/RFVZ2UT31wbCb/tJZw5zF+efZ8BWdliIVYffSZ4nz8rI81qKobHTQSpTBhrb
Rayh0qIAJ+ij15IfDkSSbCGHnccZ2pvT/VCzaZWTeGP23qjYegNpt4Vr2DephoOA4EHAB9+A3Jqi
BCe9k/VBMde3oy+74iLRP3VQmR93sIRlGDHWwv7In3KguO6sw+w8tluIxCH4GhHZzv4xghLlmRZN
UbUP0hhfyoCmUdY4EQekXkjr/Q6p1ka0GxKNDcqxo42N7YOlYgCxlYxOhVJVZR3vWh1SvkRdTfUX
ohd2lwOuNAWlLm0Kt5qrQySTDjsqPyiF36C7+AHeuaIyBJryCbTLKqZDdYRS7rX7EYbLBMqRtCmK
i2CShMaK45fguEBxhf12U5hPUwErX90oMdh4FIvnSkh0S5QhYKuMqL82sS+tbOofWbtyHqUjjtkg
GGyhKDTtLWQEEQ/Run2D/6PjMLsSo7SNubqadZgaqL6yOJV2/xA3xzJW5tMJ8kX8BAXG/n4GpGZJ
qxbAkDvbHP1N12p2/lpYx2U+do/aHIOUSjhkzX/+78/J5Z50Z/X+8mNEp9dnT1sjlukD8PUOvJca
FfTJPLENo2vEPNwfI9TPAJAqUIdmhCb3xhaMZo4wgWdexFtkOH8wLpq+MZq+IfnodTxlnYeEOtcP
31kTEBULHsDHtXH9FDubibjpQkMKXvnSQ698UuI+5xjl8uNCuP+8egiFERipCIEdw3ZbXOt0yien
nyLhUtVFUZKk7/EFNmez4ZZOfJRxVmGHSebyyU5uAyrxE5oWOzQQkJfgIkjJyidrk2WcqnX3LzVY
1HgvYC8TG6OFZjzfCAO7wL9xU3LgiqqSr9shc7gApcjBckyuzwfxyBK5V1A4eFaae+O8bNeVzHPR
CJhVCGARxK/S2pJ57KdG/ukmjHDG6YQuibePs44notHRd6mle0+wFe2uBx+DG4im4K6KKf7z4h65
w58Tyi7+eG0WR1uik5e2p/i8gsf1dPLfajBIW5AplS3bnlOOYaquURCAFlIQ9b1tMfjX5eOn1yLB
VHn0Cp2qCFepEQT5B03ua7r2X8+YNfmtEdxvcdSts8CN3FEfxoOZklH5AFSunDKJNGz2oHkclhJG
2rN7XirY3fUbO/rkOvpiT97cMIwbkHts0whOPHhuSQbGsORYwD/sW/qFzSY7jl7SWiLt+RCwmHET
IcS+bVNOH/Mfko3OC3nDaYDuKYzbsCjBw8hm43juJfcV5m9BiZ9Locms+qVagMhpbJGM6nJl2fwy
X1RuprjY+M50+Ohk8F7tTQIlRjgIkTpsZd6fVH/SGI01PFiZOjA2Zo7ic2W65jIpyChMJytfIW+Q
BntxeUjUeh2lMmmFllDuQfgURZ/YH00ZEyuRm7YmZV1HmaiDIyw3v7pa8AcnQ19t/wFB9E2t3/an
IZgI3WJu8CLYEUD6/2SXhTZlrlpAWRntOvw5O320Vvxf5tWC0uYJtsvvZptkbSDMii5JFBQm0RM2
RMcIboCX+w5N0dmAK45p1cuUokzInKDIMit6saWOv0fDiPs2RdT2YTaBw7jHYjeJgUvc2+loQ09g
gbkD6ekfcWpb9/hIzyvozpTvdue2hBBOlUEae0Logyp8rE74gRR4ephMsd3GEGOdNHJwbjT44rs9
EaEY0VCc3xSF3gyPAYbQRgN/UyV1IojYfjLi7EbraqcsmRMphWTus8j6ob+l55JZYMHRYErRW09i
NelmHjrGlcB1Sp4N/NTCeV/ng5igevkVxGXnyaHbiprcrHGQtDjmsn/p9aZ4RTGXzhdthf6FsOhh
i5PTkidsWHT7J0s7t4GNbDS1fD5SHG+ygUkqB92XfHgWID29N7/xCxkNLin/OVNE3uTqP08H2NqK
LXTmroOxNM2AZtjNvTqa+AWZkvMAE8oe7iam9gkGo7ZSD0sb8pyA46Vbi7L2jCuj9f9JLbvlAARZ
Fy/bezU5hpCquy6PlZYApdwtMWd4igXedFndaRHdDy6+fGK50s09vCs1U5hG517u48WxU9i+M4iV
eG61IJNec0GNj0A=
`protect end_protected
